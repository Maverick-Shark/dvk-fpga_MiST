library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c4f9c287",
    12 => x"86c0c64e",
    13 => x"49c4f9c2",
    14 => x"48d0e6c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087cae0",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48111e4f",
    50 => x"7808d4ff",
    51 => x"c14866c4",
    52 => x"58a6c888",
    53 => x"ed059870",
    54 => x"1e4f2687",
    55 => x"c348d4ff",
    56 => x"516878ff",
    57 => x"c14866c4",
    58 => x"58a6c888",
    59 => x"eb059870",
    60 => x"1e4f2687",
    61 => x"d4ff1e73",
    62 => x"7bffc34b",
    63 => x"ffc34a6b",
    64 => x"c8496b7b",
    65 => x"c3b17232",
    66 => x"4a6b7bff",
    67 => x"b27131c8",
    68 => x"6b7bffc3",
    69 => x"7232c849",
    70 => x"c44871b1",
    71 => x"264d2687",
    72 => x"264b264c",
    73 => x"5b5e0e4f",
    74 => x"710e5d5c",
    75 => x"4cd4ff4a",
    76 => x"ffc34972",
    77 => x"c27c7199",
    78 => x"05bfd0e6",
    79 => x"66d087c8",
    80 => x"d430c948",
    81 => x"66d058a6",
    82 => x"c329d849",
    83 => x"7c7199ff",
    84 => x"d04966d0",
    85 => x"99ffc329",
    86 => x"66d07c71",
    87 => x"c329c849",
    88 => x"7c7199ff",
    89 => x"c34966d0",
    90 => x"7c7199ff",
    91 => x"29d04972",
    92 => x"7199ffc3",
    93 => x"c94b6c7c",
    94 => x"c34dfff0",
    95 => x"d005abff",
    96 => x"7cffc387",
    97 => x"8dc14b6c",
    98 => x"c387c602",
    99 => x"f002abff",
   100 => x"fe487387",
   101 => x"c01e87c7",
   102 => x"48d4ff49",
   103 => x"c178ffc3",
   104 => x"b7c8c381",
   105 => x"87f104a9",
   106 => x"731e4f26",
   107 => x"c487e71e",
   108 => x"c04bdff8",
   109 => x"f0ffc01e",
   110 => x"fd49f7c1",
   111 => x"86c487e7",
   112 => x"c005a8c1",
   113 => x"d4ff87ea",
   114 => x"78ffc348",
   115 => x"c0c0c0c1",
   116 => x"c01ec0c0",
   117 => x"e9c1f0e1",
   118 => x"87c9fd49",
   119 => x"987086c4",
   120 => x"ff87ca05",
   121 => x"ffc348d4",
   122 => x"cb48c178",
   123 => x"87e6fe87",
   124 => x"fe058bc1",
   125 => x"48c087fd",
   126 => x"1e87e6fc",
   127 => x"d4ff1e73",
   128 => x"78ffc348",
   129 => x"1ec04bd3",
   130 => x"c1f0ffc0",
   131 => x"d4fc49c1",
   132 => x"7086c487",
   133 => x"87ca0598",
   134 => x"c348d4ff",
   135 => x"48c178ff",
   136 => x"f1fd87cb",
   137 => x"058bc187",
   138 => x"c087dbff",
   139 => x"87f1fb48",
   140 => x"5c5b5e0e",
   141 => x"4cd4ff0e",
   142 => x"c687dbfd",
   143 => x"e1c01eea",
   144 => x"49c8c1f0",
   145 => x"c487defb",
   146 => x"02a8c186",
   147 => x"eafe87c8",
   148 => x"c148c087",
   149 => x"dafa87e2",
   150 => x"cf497087",
   151 => x"c699ffff",
   152 => x"c802a9ea",
   153 => x"87d3fe87",
   154 => x"cbc148c0",
   155 => x"7cffc387",
   156 => x"fc4bf1c0",
   157 => x"987087f4",
   158 => x"87ebc002",
   159 => x"ffc01ec0",
   160 => x"49fac1f0",
   161 => x"c487defa",
   162 => x"05987086",
   163 => x"ffc387d9",
   164 => x"c3496c7c",
   165 => x"7c7c7cff",
   166 => x"99c0c17c",
   167 => x"c187c402",
   168 => x"c087d548",
   169 => x"c287d148",
   170 => x"87c405ab",
   171 => x"87c848c0",
   172 => x"fe058bc1",
   173 => x"48c087fd",
   174 => x"1e87e4f9",
   175 => x"e6c21e73",
   176 => x"78c148d0",
   177 => x"d0ff4bc7",
   178 => x"fb78c248",
   179 => x"d0ff87c8",
   180 => x"c078c348",
   181 => x"d0e5c01e",
   182 => x"f949c0c1",
   183 => x"86c487c7",
   184 => x"c105a8c1",
   185 => x"abc24b87",
   186 => x"c087c505",
   187 => x"87f9c048",
   188 => x"ff058bc1",
   189 => x"f7fc87d0",
   190 => x"d4e6c287",
   191 => x"05987058",
   192 => x"1ec187cd",
   193 => x"c1f0ffc0",
   194 => x"d8f849d0",
   195 => x"ff86c487",
   196 => x"ffc348d4",
   197 => x"87e0c478",
   198 => x"58d8e6c2",
   199 => x"c248d0ff",
   200 => x"48d4ff78",
   201 => x"c178ffc3",
   202 => x"87f5f748",
   203 => x"5c5b5e0e",
   204 => x"4a710e5d",
   205 => x"ff4dffc3",
   206 => x"7c754cd4",
   207 => x"c448d0ff",
   208 => x"7c7578c3",
   209 => x"ffc01e72",
   210 => x"49d8c1f0",
   211 => x"c487d6f7",
   212 => x"02987086",
   213 => x"48c087c5",
   214 => x"7587f0c0",
   215 => x"7cfec37c",
   216 => x"d41ec0c8",
   217 => x"dcf54966",
   218 => x"7586c487",
   219 => x"757c757c",
   220 => x"e0dad87c",
   221 => x"6c7c754b",
   222 => x"c5059949",
   223 => x"058bc187",
   224 => x"7c7587f3",
   225 => x"c248d0ff",
   226 => x"f648c178",
   227 => x"ff1e87cf",
   228 => x"d0ff4ad4",
   229 => x"78d1c448",
   230 => x"c17affc3",
   231 => x"87f80589",
   232 => x"731e4f26",
   233 => x"c54b711e",
   234 => x"4adfcdee",
   235 => x"c348d4ff",
   236 => x"486878ff",
   237 => x"02a8fec3",
   238 => x"8ac187c5",
   239 => x"7287ed05",
   240 => x"87c5059a",
   241 => x"eac048c0",
   242 => x"029b7387",
   243 => x"66c887cc",
   244 => x"f449731e",
   245 => x"86c487c5",
   246 => x"66c887c6",
   247 => x"87eefe49",
   248 => x"c348d4ff",
   249 => x"737878ff",
   250 => x"87c5059b",
   251 => x"d048d0ff",
   252 => x"f448c178",
   253 => x"731e87eb",
   254 => x"c04a711e",
   255 => x"48d4ff4b",
   256 => x"ff78ffc3",
   257 => x"c3c448d0",
   258 => x"48d4ff78",
   259 => x"7278ffc3",
   260 => x"f0ffc01e",
   261 => x"f449d1c1",
   262 => x"86c487cb",
   263 => x"cd059870",
   264 => x"1ec0c887",
   265 => x"fd4966cc",
   266 => x"86c487f8",
   267 => x"d0ff4b70",
   268 => x"7378c248",
   269 => x"87e9f348",
   270 => x"5c5b5e0e",
   271 => x"1ec00e5d",
   272 => x"c1f0ffc0",
   273 => x"dcf349c9",
   274 => x"c21ed287",
   275 => x"fd49d8e6",
   276 => x"86c887d0",
   277 => x"84c14cc0",
   278 => x"04acb7d2",
   279 => x"e6c287f8",
   280 => x"49bf97d8",
   281 => x"c199c0c3",
   282 => x"c005a9c0",
   283 => x"e6c287e7",
   284 => x"49bf97df",
   285 => x"e6c231d0",
   286 => x"4abf97e0",
   287 => x"b17232c8",
   288 => x"97e1e6c2",
   289 => x"71b14abf",
   290 => x"ffffcf4c",
   291 => x"84c19cff",
   292 => x"e7c134ca",
   293 => x"e1e6c287",
   294 => x"c149bf97",
   295 => x"c299c631",
   296 => x"bf97e2e6",
   297 => x"2ab7c74a",
   298 => x"e6c2b172",
   299 => x"4abf97dd",
   300 => x"c29dcf4d",
   301 => x"bf97dee6",
   302 => x"ca9ac34a",
   303 => x"dfe6c232",
   304 => x"c24bbf97",
   305 => x"c2b27333",
   306 => x"bf97e0e6",
   307 => x"9bc0c34b",
   308 => x"732bb7c6",
   309 => x"c181c2b2",
   310 => x"70307148",
   311 => x"7548c149",
   312 => x"724d7030",
   313 => x"7184c14c",
   314 => x"b7c0c894",
   315 => x"87cc06ad",
   316 => x"2db734c1",
   317 => x"adb7c0c8",
   318 => x"87f4ff01",
   319 => x"dcf04874",
   320 => x"5b5e0e87",
   321 => x"f80e5d5c",
   322 => x"feeec286",
   323 => x"c278c048",
   324 => x"c01ef6e6",
   325 => x"87defb49",
   326 => x"987086c4",
   327 => x"c087c505",
   328 => x"87cec948",
   329 => x"7ec14dc0",
   330 => x"bfcbf2c0",
   331 => x"ece7c249",
   332 => x"4bc8714a",
   333 => x"7087f3ec",
   334 => x"87c20598",
   335 => x"f2c07ec0",
   336 => x"c249bfc7",
   337 => x"714ac8e8",
   338 => x"ddec4bc8",
   339 => x"05987087",
   340 => x"7ec087c2",
   341 => x"fdc0026e",
   342 => x"fcedc287",
   343 => x"eec24dbf",
   344 => x"7ebf9ff4",
   345 => x"ead6c548",
   346 => x"87c705a8",
   347 => x"bffcedc2",
   348 => x"6e87ce4d",
   349 => x"d5e9ca48",
   350 => x"87c502a8",
   351 => x"f1c748c0",
   352 => x"f6e6c287",
   353 => x"f949751e",
   354 => x"86c487ec",
   355 => x"c5059870",
   356 => x"c748c087",
   357 => x"f2c087dc",
   358 => x"c249bfc7",
   359 => x"714ac8e8",
   360 => x"c5eb4bc8",
   361 => x"05987087",
   362 => x"eec287c8",
   363 => x"78c148fe",
   364 => x"f2c087da",
   365 => x"c249bfcb",
   366 => x"714aece7",
   367 => x"e9ea4bc8",
   368 => x"02987087",
   369 => x"c087c5c0",
   370 => x"87e6c648",
   371 => x"97f4eec2",
   372 => x"d5c149bf",
   373 => x"cdc005a9",
   374 => x"f5eec287",
   375 => x"c249bf97",
   376 => x"c002a9ea",
   377 => x"48c087c5",
   378 => x"c287c7c6",
   379 => x"bf97f6e6",
   380 => x"e9c3487e",
   381 => x"cec002a8",
   382 => x"c3486e87",
   383 => x"c002a8eb",
   384 => x"48c087c5",
   385 => x"c287ebc5",
   386 => x"bf97c1e7",
   387 => x"c0059949",
   388 => x"e7c287cc",
   389 => x"49bf97c2",
   390 => x"c002a9c2",
   391 => x"48c087c5",
   392 => x"c287cfc5",
   393 => x"bf97c3e7",
   394 => x"faeec248",
   395 => x"484c7058",
   396 => x"eec288c1",
   397 => x"e7c258fe",
   398 => x"49bf97c4",
   399 => x"e7c28175",
   400 => x"4abf97c5",
   401 => x"a17232c8",
   402 => x"cbf3c27e",
   403 => x"c2786e48",
   404 => x"bf97c6e7",
   405 => x"58a6c848",
   406 => x"bffeeec2",
   407 => x"87d4c202",
   408 => x"bfc7f2c0",
   409 => x"c8e8c249",
   410 => x"4bc8714a",
   411 => x"7087fbe7",
   412 => x"c5c00298",
   413 => x"c348c087",
   414 => x"eec287f8",
   415 => x"c24cbff6",
   416 => x"c25cdff3",
   417 => x"bf97dbe7",
   418 => x"c231c849",
   419 => x"bf97dae7",
   420 => x"c249a14a",
   421 => x"bf97dce7",
   422 => x"7232d04a",
   423 => x"e7c249a1",
   424 => x"4abf97dd",
   425 => x"a17232d8",
   426 => x"9166c449",
   427 => x"bfcbf3c2",
   428 => x"d3f3c281",
   429 => x"e3e7c259",
   430 => x"c84abf97",
   431 => x"e2e7c232",
   432 => x"a24bbf97",
   433 => x"e4e7c24a",
   434 => x"d04bbf97",
   435 => x"4aa27333",
   436 => x"97e5e7c2",
   437 => x"9bcf4bbf",
   438 => x"a27333d8",
   439 => x"d7f3c24a",
   440 => x"d3f3c25a",
   441 => x"8ac24abf",
   442 => x"f3c29274",
   443 => x"a17248d7",
   444 => x"87cac178",
   445 => x"97c8e7c2",
   446 => x"31c849bf",
   447 => x"97c7e7c2",
   448 => x"49a14abf",
   449 => x"59c6efc2",
   450 => x"bfc2efc2",
   451 => x"c731c549",
   452 => x"29c981ff",
   453 => x"59dff3c2",
   454 => x"97cde7c2",
   455 => x"32c84abf",
   456 => x"97cce7c2",
   457 => x"4aa24bbf",
   458 => x"6e9266c4",
   459 => x"dbf3c282",
   460 => x"d3f3c25a",
   461 => x"c278c048",
   462 => x"7248cff3",
   463 => x"f3c278a1",
   464 => x"f3c248df",
   465 => x"c278bfd3",
   466 => x"c248e3f3",
   467 => x"78bfd7f3",
   468 => x"bffeeec2",
   469 => x"87c9c002",
   470 => x"30c44874",
   471 => x"c9c07e70",
   472 => x"dbf3c287",
   473 => x"30c448bf",
   474 => x"efc27e70",
   475 => x"786e48c2",
   476 => x"8ef848c1",
   477 => x"4c264d26",
   478 => x"4f264b26",
   479 => x"5c5b5e0e",
   480 => x"4a710e5d",
   481 => x"bffeeec2",
   482 => x"7287cb02",
   483 => x"722bc74b",
   484 => x"9cffc14c",
   485 => x"4b7287c9",
   486 => x"4c722bc8",
   487 => x"c29cffc3",
   488 => x"83bfcbf3",
   489 => x"bfc3f2c0",
   490 => x"87d902ab",
   491 => x"5bc7f2c0",
   492 => x"1ef6e6c2",
   493 => x"fdf04973",
   494 => x"7086c487",
   495 => x"87c50598",
   496 => x"e6c048c0",
   497 => x"feeec287",
   498 => x"87d202bf",
   499 => x"91c44974",
   500 => x"81f6e6c2",
   501 => x"ffcf4d69",
   502 => x"9dffffff",
   503 => x"497487cb",
   504 => x"e6c291c2",
   505 => x"699f81f6",
   506 => x"fe48754d",
   507 => x"5e0e87c6",
   508 => x"0e5d5c5b",
   509 => x"c04d711e",
   510 => x"ca49c11e",
   511 => x"86c487ee",
   512 => x"029c4c70",
   513 => x"c287c0c1",
   514 => x"754ac6ef",
   515 => x"87ffe049",
   516 => x"c0029870",
   517 => x"4a7487f1",
   518 => x"4bcb4975",
   519 => x"7087e5e1",
   520 => x"e2c00298",
   521 => x"741ec087",
   522 => x"87c7029c",
   523 => x"c048a6c4",
   524 => x"c487c578",
   525 => x"78c148a6",
   526 => x"c94966c4",
   527 => x"86c487ee",
   528 => x"059c4c70",
   529 => x"7487c0ff",
   530 => x"e7fc2648",
   531 => x"5b5e0e87",
   532 => x"1e0e5d5c",
   533 => x"059b4b71",
   534 => x"48c087c5",
   535 => x"c887e5c1",
   536 => x"7dc04da3",
   537 => x"c70266d4",
   538 => x"9766d487",
   539 => x"87c505bf",
   540 => x"cfc148c0",
   541 => x"4966d487",
   542 => x"7087f3fd",
   543 => x"c1029c4c",
   544 => x"a4dc87c0",
   545 => x"da7d6949",
   546 => x"a3c449a4",
   547 => x"7a699f4a",
   548 => x"bffeeec2",
   549 => x"d487d202",
   550 => x"699f49a4",
   551 => x"ffffc049",
   552 => x"d0487199",
   553 => x"c27e7030",
   554 => x"6e7ec087",
   555 => x"806a4849",
   556 => x"7bc07a70",
   557 => x"6a49a3cc",
   558 => x"49a3d079",
   559 => x"487479c0",
   560 => x"48c087c2",
   561 => x"87ecfa26",
   562 => x"5c5b5e0e",
   563 => x"4c710e5d",
   564 => x"48c3f2c0",
   565 => x"9c7478ff",
   566 => x"87cac102",
   567 => x"6949a4c8",
   568 => x"87c2c102",
   569 => x"6c4a66d0",
   570 => x"a6d48249",
   571 => x"4d66d05a",
   572 => x"faeec2b9",
   573 => x"baff4abf",
   574 => x"99719972",
   575 => x"87e4c002",
   576 => x"6b4ba4c4",
   577 => x"87f4f949",
   578 => x"eec27b70",
   579 => x"6c49bff6",
   580 => x"757c7181",
   581 => x"faeec2b9",
   582 => x"baff4abf",
   583 => x"99719972",
   584 => x"87dcff05",
   585 => x"cbf97c75",
   586 => x"1e731e87",
   587 => x"029b4b71",
   588 => x"a3c887c7",
   589 => x"c5056949",
   590 => x"c048c087",
   591 => x"f3c287eb",
   592 => x"c44abfcf",
   593 => x"496949a3",
   594 => x"eec289c2",
   595 => x"7191bff6",
   596 => x"eec24aa2",
   597 => x"6b49bffa",
   598 => x"4aa27199",
   599 => x"721e66c8",
   600 => x"87d2ea49",
   601 => x"497086c4",
   602 => x"87ccf848",
   603 => x"711e731e",
   604 => x"c7029b4b",
   605 => x"49a3c887",
   606 => x"87c50569",
   607 => x"ebc048c0",
   608 => x"cff3c287",
   609 => x"a3c44abf",
   610 => x"c2496949",
   611 => x"f6eec289",
   612 => x"a27191bf",
   613 => x"faeec24a",
   614 => x"996b49bf",
   615 => x"c84aa271",
   616 => x"49721e66",
   617 => x"c487c5e6",
   618 => x"48497086",
   619 => x"0e87c9f7",
   620 => x"5d5c5b5e",
   621 => x"4b711e0e",
   622 => x"c94c66d4",
   623 => x"029b732c",
   624 => x"c887cfc1",
   625 => x"026949a3",
   626 => x"d087c7c1",
   627 => x"66d44da3",
   628 => x"faeec27d",
   629 => x"b9ff49bf",
   630 => x"7e994a6b",
   631 => x"cd03ac71",
   632 => x"7d7bc087",
   633 => x"c44aa3cc",
   634 => x"796a49a3",
   635 => x"8c7287c2",
   636 => x"dd029c74",
   637 => x"731e4987",
   638 => x"87ccfb49",
   639 => x"66d486c4",
   640 => x"99ffc749",
   641 => x"c287cb02",
   642 => x"731ef6e6",
   643 => x"87d9fc49",
   644 => x"f52686c4",
   645 => x"731e87de",
   646 => x"9b4b711e",
   647 => x"87e4c002",
   648 => x"5be3f3c2",
   649 => x"8ac24a73",
   650 => x"bff6eec2",
   651 => x"f3c29249",
   652 => x"7248bfcf",
   653 => x"e7f3c280",
   654 => x"c4487158",
   655 => x"c6efc230",
   656 => x"87edc058",
   657 => x"48dff3c2",
   658 => x"bfd3f3c2",
   659 => x"e3f3c278",
   660 => x"d7f3c248",
   661 => x"eec278bf",
   662 => x"c902bffe",
   663 => x"f6eec287",
   664 => x"31c449bf",
   665 => x"f3c287c7",
   666 => x"c449bfdb",
   667 => x"c6efc231",
   668 => x"87c4f459",
   669 => x"5c5b5e0e",
   670 => x"c04a710e",
   671 => x"029a724b",
   672 => x"da87e1c0",
   673 => x"699f49a2",
   674 => x"feeec24b",
   675 => x"87cf02bf",
   676 => x"9f49a2d4",
   677 => x"c04c4969",
   678 => x"d09cffff",
   679 => x"c087c234",
   680 => x"b349744c",
   681 => x"edfd4973",
   682 => x"87caf387",
   683 => x"5c5b5e0e",
   684 => x"86f40e5d",
   685 => x"7ec04a71",
   686 => x"d8029a72",
   687 => x"f2e6c287",
   688 => x"c278c048",
   689 => x"c248eae6",
   690 => x"78bfe3f3",
   691 => x"48eee6c2",
   692 => x"bfdff3c2",
   693 => x"d3efc278",
   694 => x"c250c048",
   695 => x"49bfc2ef",
   696 => x"bff2e6c2",
   697 => x"03aa714a",
   698 => x"7287ffc3",
   699 => x"0599cf49",
   700 => x"c287e0c0",
   701 => x"c21ef6e6",
   702 => x"49bfeae6",
   703 => x"48eae6c2",
   704 => x"7178a1c1",
   705 => x"c487efe3",
   706 => x"fff1c086",
   707 => x"f6e6c248",
   708 => x"c087cc78",
   709 => x"48bffff1",
   710 => x"c080e0c0",
   711 => x"c258c3f2",
   712 => x"48bff2e6",
   713 => x"e6c280c1",
   714 => x"7f2758f6",
   715 => x"bf00000c",
   716 => x"9d4dbf97",
   717 => x"87e2c202",
   718 => x"02ade5c3",
   719 => x"c087dbc2",
   720 => x"4bbffff1",
   721 => x"1149a3cb",
   722 => x"05accf4c",
   723 => x"7587d2c1",
   724 => x"c199df49",
   725 => x"c291cd89",
   726 => x"c181c6ef",
   727 => x"51124aa3",
   728 => x"124aa3c3",
   729 => x"4aa3c551",
   730 => x"a3c75112",
   731 => x"c951124a",
   732 => x"51124aa3",
   733 => x"124aa3ce",
   734 => x"4aa3d051",
   735 => x"a3d25112",
   736 => x"d451124a",
   737 => x"51124aa3",
   738 => x"124aa3d6",
   739 => x"4aa3d851",
   740 => x"a3dc5112",
   741 => x"de51124a",
   742 => x"51124aa3",
   743 => x"f9c07ec1",
   744 => x"c8497487",
   745 => x"eac00599",
   746 => x"d0497487",
   747 => x"87d00599",
   748 => x"c00266dc",
   749 => x"497387ca",
   750 => x"700f66dc",
   751 => x"87d30298",
   752 => x"c6c0056e",
   753 => x"c6efc287",
   754 => x"c050c048",
   755 => x"48bffff1",
   756 => x"c287e7c2",
   757 => x"c048d3ef",
   758 => x"efc27e50",
   759 => x"c249bfc2",
   760 => x"4abff2e6",
   761 => x"fc04aa71",
   762 => x"f3c287c1",
   763 => x"c005bfe3",
   764 => x"eec287c8",
   765 => x"c102bffe",
   766 => x"f2c087fe",
   767 => x"78ff48c3",
   768 => x"bfeee6c2",
   769 => x"87f4ed49",
   770 => x"e6c24970",
   771 => x"a6c459f2",
   772 => x"eee6c248",
   773 => x"eec278bf",
   774 => x"c002bffe",
   775 => x"66c487d8",
   776 => x"ffffcf49",
   777 => x"a999f8ff",
   778 => x"87c5c002",
   779 => x"e1c04dc0",
   780 => x"c04dc187",
   781 => x"66c487dc",
   782 => x"f8ffcf49",
   783 => x"c002a999",
   784 => x"a6c887c8",
   785 => x"c078c048",
   786 => x"a6c887c5",
   787 => x"c878c148",
   788 => x"9d754d66",
   789 => x"87e0c005",
   790 => x"c24966c4",
   791 => x"f6eec289",
   792 => x"c2914abf",
   793 => x"4abfcff3",
   794 => x"48eae6c2",
   795 => x"c278a172",
   796 => x"c048f2e6",
   797 => x"87e3f978",
   798 => x"8ef448c0",
   799 => x"0087f5eb",
   800 => x"ff000000",
   801 => x"8fffffff",
   802 => x"9800000c",
   803 => x"4600000c",
   804 => x"32335441",
   805 => x"00202020",
   806 => x"31544146",
   807 => x"20202036",
   808 => x"d4ff1e00",
   809 => x"78ffc348",
   810 => x"4f264868",
   811 => x"48d4ff1e",
   812 => x"ff78ffc3",
   813 => x"e1c848d0",
   814 => x"48d4ff78",
   815 => x"f3c278d4",
   816 => x"d4ff48e7",
   817 => x"4f2650bf",
   818 => x"48d0ff1e",
   819 => x"2678e0c0",
   820 => x"ccff1e4f",
   821 => x"99497087",
   822 => x"c087c602",
   823 => x"f105a9fb",
   824 => x"26487187",
   825 => x"5b5e0e4f",
   826 => x"4b710e5c",
   827 => x"f0fe4cc0",
   828 => x"99497087",
   829 => x"87f9c002",
   830 => x"02a9ecc0",
   831 => x"c087f2c0",
   832 => x"c002a9fb",
   833 => x"66cc87eb",
   834 => x"c703acb7",
   835 => x"0266d087",
   836 => x"537187c2",
   837 => x"c2029971",
   838 => x"fe84c187",
   839 => x"497087c3",
   840 => x"87cd0299",
   841 => x"02a9ecc0",
   842 => x"fbc087c7",
   843 => x"d5ff05a9",
   844 => x"0266d087",
   845 => x"97c087c3",
   846 => x"a9ecc07b",
   847 => x"7487c405",
   848 => x"7487c54a",
   849 => x"8a0ac04a",
   850 => x"87c24872",
   851 => x"4c264d26",
   852 => x"4f264b26",
   853 => x"87c9fd1e",
   854 => x"f0c04970",
   855 => x"ca04a9b7",
   856 => x"b7f9c087",
   857 => x"87c301a9",
   858 => x"c189f0c0",
   859 => x"04a9b7c1",
   860 => x"dac187ca",
   861 => x"c301a9b7",
   862 => x"89f7c087",
   863 => x"4f264871",
   864 => x"5c5b5e0e",
   865 => x"ff4a710e",
   866 => x"49724cd4",
   867 => x"7087eac0",
   868 => x"c2029b4b",
   869 => x"ff8bc187",
   870 => x"c5c848d0",
   871 => x"7cd5c178",
   872 => x"31c64973",
   873 => x"97c9e3c2",
   874 => x"71484abf",
   875 => x"ff7c70b0",
   876 => x"78c448d0",
   877 => x"d5fe4873",
   878 => x"5b5e0e87",
   879 => x"f80e5d5c",
   880 => x"c04b7186",
   881 => x"e0fac07e",
   882 => x"df49bf97",
   883 => x"eec005a9",
   884 => x"49a3c887",
   885 => x"c1496997",
   886 => x"dd05a9c3",
   887 => x"49a3c987",
   888 => x"c1496997",
   889 => x"d105a9c6",
   890 => x"49a3ca87",
   891 => x"c1496997",
   892 => x"c505a9c7",
   893 => x"c248c187",
   894 => x"48c087e1",
   895 => x"fa87dcc2",
   896 => x"4cc087ea",
   897 => x"97e0fac0",
   898 => x"a9c049bf",
   899 => x"fa87cf04",
   900 => x"84c187ff",
   901 => x"97e0fac0",
   902 => x"06ac49bf",
   903 => x"fac087f1",
   904 => x"02bf97e0",
   905 => x"f8f987cf",
   906 => x"99497087",
   907 => x"c087c602",
   908 => x"f105a9ec",
   909 => x"f94cc087",
   910 => x"4d7087e7",
   911 => x"c887e2f9",
   912 => x"dcf958a6",
   913 => x"c14a7087",
   914 => x"49a3c884",
   915 => x"ad496997",
   916 => x"c087c702",
   917 => x"c005adff",
   918 => x"a3c987e7",
   919 => x"49699749",
   920 => x"02a966c4",
   921 => x"c04887c7",
   922 => x"d405a8ff",
   923 => x"49a3ca87",
   924 => x"aa496997",
   925 => x"c087c602",
   926 => x"c405aaff",
   927 => x"d07ec187",
   928 => x"adecc087",
   929 => x"c087c602",
   930 => x"c405adfb",
   931 => x"c14cc087",
   932 => x"fe026e7e",
   933 => x"eff887e1",
   934 => x"f8487487",
   935 => x"87ecfa8e",
   936 => x"5b5e0e00",
   937 => x"1e0e5d5c",
   938 => x"4cc04b71",
   939 => x"c004ab4d",
   940 => x"f6c087e8",
   941 => x"9d751ef9",
   942 => x"c087c402",
   943 => x"c187c24a",
   944 => x"ef49724a",
   945 => x"86c487e6",
   946 => x"84c17e70",
   947 => x"87c2056e",
   948 => x"85c14c73",
   949 => x"ff06ac73",
   950 => x"486e87d8",
   951 => x"264d2626",
   952 => x"264b264c",
   953 => x"5b5e0e4f",
   954 => x"1e0e5d5c",
   955 => x"de494c71",
   956 => x"c1f4c291",
   957 => x"9785714d",
   958 => x"ddc1026d",
   959 => x"ecf3c287",
   960 => x"82744abf",
   961 => x"d8fe4972",
   962 => x"6e7e7087",
   963 => x"87f3c002",
   964 => x"4bf4f3c2",
   965 => x"49cb4a6e",
   966 => x"87ccc6ff",
   967 => x"93cb4b74",
   968 => x"83dce2c1",
   969 => x"fdc083c4",
   970 => x"49747bde",
   971 => x"87d6c7c1",
   972 => x"f4c27b75",
   973 => x"49bf97c0",
   974 => x"f4f3c21e",
   975 => x"ece4c149",
   976 => x"7486c487",
   977 => x"fdc6c149",
   978 => x"c149c087",
   979 => x"c287dcc8",
   980 => x"c048e8f3",
   981 => x"df49c178",
   982 => x"fd2687fd",
   983 => x"6f4c87ff",
   984 => x"6e696461",
   985 => x"2e2e2e67",
   986 => x"5b5e0e00",
   987 => x"4b710e5c",
   988 => x"ecf3c24a",
   989 => x"497282bf",
   990 => x"7087e6fc",
   991 => x"c4029c4c",
   992 => x"efeb4987",
   993 => x"ecf3c287",
   994 => x"c178c048",
   995 => x"87c7df49",
   996 => x"0e87ccfd",
   997 => x"5d5c5b5e",
   998 => x"c286f40e",
   999 => x"c04df6e6",
  1000 => x"48a6c44c",
  1001 => x"f3c278c0",
  1002 => x"c049bfec",
  1003 => x"c1c106a9",
  1004 => x"f6e6c287",
  1005 => x"c0029848",
  1006 => x"f6c087f8",
  1007 => x"66c81ef9",
  1008 => x"c487c702",
  1009 => x"78c048a6",
  1010 => x"a6c487c5",
  1011 => x"c478c148",
  1012 => x"d7eb4966",
  1013 => x"7086c487",
  1014 => x"c484c14d",
  1015 => x"80c14866",
  1016 => x"c258a6c8",
  1017 => x"49bfecf3",
  1018 => x"87c603ac",
  1019 => x"ff059d75",
  1020 => x"4cc087c8",
  1021 => x"c3029d75",
  1022 => x"f6c087e0",
  1023 => x"66c81ef9",
  1024 => x"cc87c702",
  1025 => x"78c048a6",
  1026 => x"a6cc87c5",
  1027 => x"cc78c148",
  1028 => x"d7ea4966",
  1029 => x"7086c487",
  1030 => x"c2026e7e",
  1031 => x"496e87e9",
  1032 => x"699781cb",
  1033 => x"0299d049",
  1034 => x"c087d6c1",
  1035 => x"744ae9fd",
  1036 => x"c191cb49",
  1037 => x"7281dce2",
  1038 => x"c381c879",
  1039 => x"497451ff",
  1040 => x"f4c291de",
  1041 => x"85714dc1",
  1042 => x"7d97c1c2",
  1043 => x"c049a5c1",
  1044 => x"efc251e0",
  1045 => x"02bf97c6",
  1046 => x"84c187d2",
  1047 => x"c24ba5c2",
  1048 => x"db4ac6ef",
  1049 => x"ffc0ff49",
  1050 => x"87dbc187",
  1051 => x"c049a5cd",
  1052 => x"c284c151",
  1053 => x"4a6e4ba5",
  1054 => x"c0ff49cb",
  1055 => x"c6c187ea",
  1056 => x"e5fbc087",
  1057 => x"cb49744a",
  1058 => x"dce2c191",
  1059 => x"c2797281",
  1060 => x"bf97c6ef",
  1061 => x"7487d802",
  1062 => x"c191de49",
  1063 => x"c1f4c284",
  1064 => x"c283714b",
  1065 => x"dd4ac6ef",
  1066 => x"fbfffe49",
  1067 => x"7487d887",
  1068 => x"c293de4b",
  1069 => x"cb83c1f4",
  1070 => x"51c049a3",
  1071 => x"6e7384c1",
  1072 => x"fe49cb4a",
  1073 => x"c487e1ff",
  1074 => x"80c14866",
  1075 => x"c758a6c8",
  1076 => x"c5c003ac",
  1077 => x"fc056e87",
  1078 => x"487487e0",
  1079 => x"fcf78ef4",
  1080 => x"1e731e87",
  1081 => x"cb494b71",
  1082 => x"dce2c191",
  1083 => x"4aa1c881",
  1084 => x"48c9e3c2",
  1085 => x"a1c95012",
  1086 => x"e0fac04a",
  1087 => x"ca501248",
  1088 => x"c0f4c281",
  1089 => x"c2501148",
  1090 => x"bf97c0f4",
  1091 => x"49c01e49",
  1092 => x"87d9ddc1",
  1093 => x"48e8f3c2",
  1094 => x"49c178de",
  1095 => x"2687f8d8",
  1096 => x"1e87fef6",
  1097 => x"cb494a71",
  1098 => x"dce2c191",
  1099 => x"1181c881",
  1100 => x"ecf3c248",
  1101 => x"ecf3c258",
  1102 => x"c178c048",
  1103 => x"87d7d849",
  1104 => x"c01e4f26",
  1105 => x"e2c0c149",
  1106 => x"1e4f2687",
  1107 => x"d2029971",
  1108 => x"f1e3c187",
  1109 => x"f750c048",
  1110 => x"e3c4c180",
  1111 => x"cae2c140",
  1112 => x"c187ce78",
  1113 => x"c148ede3",
  1114 => x"fc78ebe1",
  1115 => x"c2c5c180",
  1116 => x"0e4f2678",
  1117 => x"0e5c5b5e",
  1118 => x"cb4a4c71",
  1119 => x"dce2c192",
  1120 => x"49a2c882",
  1121 => x"974ba2c9",
  1122 => x"971e4b6b",
  1123 => x"ca1e4969",
  1124 => x"c0491282",
  1125 => x"c087ddeb",
  1126 => x"87fbd649",
  1127 => x"fdc04974",
  1128 => x"8ef887e4",
  1129 => x"1e87f8f4",
  1130 => x"4b711e73",
  1131 => x"87c3ff49",
  1132 => x"fefe4973",
  1133 => x"87e9f487",
  1134 => x"711e731e",
  1135 => x"4aa3c64b",
  1136 => x"c187dc02",
  1137 => x"e4c0028a",
  1138 => x"c1028a87",
  1139 => x"028a87e8",
  1140 => x"8a87cac1",
  1141 => x"87efc002",
  1142 => x"87d9028a",
  1143 => x"c287e9c1",
  1144 => x"df48e8f3",
  1145 => x"d549c178",
  1146 => x"e6c187ed",
  1147 => x"fc49c787",
  1148 => x"dec187f1",
  1149 => x"ecf3c287",
  1150 => x"cbc102bf",
  1151 => x"88c14887",
  1152 => x"58f0f3c2",
  1153 => x"c287c1c1",
  1154 => x"02bff0f3",
  1155 => x"c287f9c0",
  1156 => x"48bfecf3",
  1157 => x"f3c280c1",
  1158 => x"ebc058f0",
  1159 => x"ecf3c287",
  1160 => x"89c649bf",
  1161 => x"59f0f3c2",
  1162 => x"03a9b7c0",
  1163 => x"f3c287da",
  1164 => x"78c048ec",
  1165 => x"f3c287d2",
  1166 => x"cb02bff0",
  1167 => x"ecf3c287",
  1168 => x"80c648bf",
  1169 => x"58f0f3c2",
  1170 => x"cad449c0",
  1171 => x"c0497387",
  1172 => x"f287f3fa",
  1173 => x"5e0e87cb",
  1174 => x"710e5c5b",
  1175 => x"1e66cc4c",
  1176 => x"93cb4b74",
  1177 => x"83dce2c1",
  1178 => x"6a4aa3c4",
  1179 => x"c7f9fe49",
  1180 => x"e1c3c187",
  1181 => x"49a3c87b",
  1182 => x"c95166d4",
  1183 => x"66d849a3",
  1184 => x"49a3ca51",
  1185 => x"265166dc",
  1186 => x"0e87d4f1",
  1187 => x"5d5c5b5e",
  1188 => x"86d0ff0e",
  1189 => x"c859a6d8",
  1190 => x"78c048a6",
  1191 => x"c4c180fc",
  1192 => x"80c87866",
  1193 => x"80c478c1",
  1194 => x"f3c278c1",
  1195 => x"78c148f0",
  1196 => x"bfe8f3c2",
  1197 => x"de486e7e",
  1198 => x"87cb05a8",
  1199 => x"7087d4f3",
  1200 => x"59a6cc49",
  1201 => x"6e87f8d0",
  1202 => x"05a8df48",
  1203 => x"c187eec1",
  1204 => x"c44966c0",
  1205 => x"c17e6981",
  1206 => x"6e48f4dc",
  1207 => x"4aa1d049",
  1208 => x"aa714120",
  1209 => x"c187f905",
  1210 => x"c14ae1c3",
  1211 => x"7a0a66c0",
  1212 => x"66c0c10a",
  1213 => x"df81c949",
  1214 => x"66c0c151",
  1215 => x"c181ca49",
  1216 => x"c0c151d3",
  1217 => x"81cb4966",
  1218 => x"c44ba1c4",
  1219 => x"786b48a6",
  1220 => x"1e721e71",
  1221 => x"48c4ddc1",
  1222 => x"d04966cc",
  1223 => x"41204aa1",
  1224 => x"f905aa71",
  1225 => x"264a2687",
  1226 => x"c9797249",
  1227 => x"52df4aa1",
  1228 => x"d4c181ca",
  1229 => x"48a6c851",
  1230 => x"c2cf78c2",
  1231 => x"87ece587",
  1232 => x"e587cee6",
  1233 => x"4c7087db",
  1234 => x"02acfbc0",
  1235 => x"d487d0c1",
  1236 => x"c2c10566",
  1237 => x"1e1ec087",
  1238 => x"e4c11ec1",
  1239 => x"49c01ed2",
  1240 => x"c187f3fb",
  1241 => x"c44a66d0",
  1242 => x"c7496a82",
  1243 => x"c1517481",
  1244 => x"6a1ed81e",
  1245 => x"e581c849",
  1246 => x"86d887eb",
  1247 => x"4866c4c1",
  1248 => x"c701a8c0",
  1249 => x"48a6c887",
  1250 => x"87ce78c1",
  1251 => x"4866c4c1",
  1252 => x"a6c888c1",
  1253 => x"e487c358",
  1254 => x"a6cc87f7",
  1255 => x"7478c248",
  1256 => x"d6cd029c",
  1257 => x"4866c887",
  1258 => x"a866c8c1",
  1259 => x"87cbcd03",
  1260 => x"c048a6d8",
  1261 => x"87e9e378",
  1262 => x"d0c14c70",
  1263 => x"d6c205ac",
  1264 => x"7e66d887",
  1265 => x"7087cde6",
  1266 => x"59a6dc49",
  1267 => x"7087d2e3",
  1268 => x"acecc04c",
  1269 => x"87eac105",
  1270 => x"cb4966c8",
  1271 => x"66c0c191",
  1272 => x"4aa1c481",
  1273 => x"a1c84d6a",
  1274 => x"5266d84a",
  1275 => x"79e3c4c1",
  1276 => x"7087eee2",
  1277 => x"d8029c4c",
  1278 => x"acfbc087",
  1279 => x"7487d202",
  1280 => x"87dde255",
  1281 => x"029c4c70",
  1282 => x"fbc087c7",
  1283 => x"eeff05ac",
  1284 => x"55e0c087",
  1285 => x"c055c1c2",
  1286 => x"66d47d97",
  1287 => x"05a96e49",
  1288 => x"66c887db",
  1289 => x"a866c448",
  1290 => x"c887ca04",
  1291 => x"80c14866",
  1292 => x"c858a6cc",
  1293 => x"4866c487",
  1294 => x"a6c888c1",
  1295 => x"87e1e158",
  1296 => x"d0c14c70",
  1297 => x"87c805ac",
  1298 => x"c14866d0",
  1299 => x"58a6d480",
  1300 => x"02acd0c1",
  1301 => x"dc87eafd",
  1302 => x"66d448a6",
  1303 => x"4866d878",
  1304 => x"05a866dc",
  1305 => x"c087e6c9",
  1306 => x"c048a6e0",
  1307 => x"80c478f0",
  1308 => x"c47866cc",
  1309 => x"7e78c080",
  1310 => x"fbc04874",
  1311 => x"a6f0c088",
  1312 => x"02987058",
  1313 => x"4887e1c8",
  1314 => x"f0c088cb",
  1315 => x"987058a6",
  1316 => x"87e9c002",
  1317 => x"c088c948",
  1318 => x"7058a6f0",
  1319 => x"e9c30298",
  1320 => x"88c44887",
  1321 => x"58a6f0c0",
  1322 => x"d6029870",
  1323 => x"88c14887",
  1324 => x"58a6f0c0",
  1325 => x"c3029870",
  1326 => x"e5c787d0",
  1327 => x"a6e0c087",
  1328 => x"cc78c048",
  1329 => x"80c14866",
  1330 => x"ff58a6d0",
  1331 => x"7087d2df",
  1332 => x"acecc04c",
  1333 => x"c087d702",
  1334 => x"c00266e0",
  1335 => x"e4c087c7",
  1336 => x"c9c05ca6",
  1337 => x"c0487487",
  1338 => x"e8c088f0",
  1339 => x"ecc058a6",
  1340 => x"cdc002ac",
  1341 => x"e8deff87",
  1342 => x"c04c7087",
  1343 => x"ff05acec",
  1344 => x"e0c087f3",
  1345 => x"66d41e66",
  1346 => x"ecc01e49",
  1347 => x"e4c11e66",
  1348 => x"66d81ed2",
  1349 => x"87fef449",
  1350 => x"1eca1ec0",
  1351 => x"4966e0c0",
  1352 => x"d8c191cb",
  1353 => x"a6d88166",
  1354 => x"78a1c448",
  1355 => x"49bf66d8",
  1356 => x"87f1deff",
  1357 => x"b7c086d8",
  1358 => x"c8c106a8",
  1359 => x"de1ec187",
  1360 => x"bf66c81e",
  1361 => x"dcdeff49",
  1362 => x"7086c887",
  1363 => x"08c04849",
  1364 => x"a6e4c088",
  1365 => x"a8b7c058",
  1366 => x"87e9c006",
  1367 => x"4866e0c0",
  1368 => x"03a8b7dd",
  1369 => x"bf6e87df",
  1370 => x"66e0c049",
  1371 => x"51e0c081",
  1372 => x"81c14966",
  1373 => x"c281bf6e",
  1374 => x"e0c051c1",
  1375 => x"81c24966",
  1376 => x"c081bf6e",
  1377 => x"c47ec151",
  1378 => x"dfff87de",
  1379 => x"e4c087c6",
  1380 => x"deff58a6",
  1381 => x"e8c087fe",
  1382 => x"ecc058a6",
  1383 => x"cbc005a8",
  1384 => x"a6e4c087",
  1385 => x"66e0c048",
  1386 => x"87c4c078",
  1387 => x"87f1dbff",
  1388 => x"cb4966c8",
  1389 => x"66c0c191",
  1390 => x"70807148",
  1391 => x"c84a6e7e",
  1392 => x"ca496e82",
  1393 => x"66e0c081",
  1394 => x"66e4c051",
  1395 => x"c081c149",
  1396 => x"c18966e0",
  1397 => x"70307148",
  1398 => x"7189c149",
  1399 => x"f7c27a97",
  1400 => x"c049bfdd",
  1401 => x"972966e0",
  1402 => x"71484a6a",
  1403 => x"a6f0c098",
  1404 => x"c4496e58",
  1405 => x"dc4d6981",
  1406 => x"66d84866",
  1407 => x"c8c002a8",
  1408 => x"48a6d887",
  1409 => x"c5c078c0",
  1410 => x"48a6d887",
  1411 => x"66d878c1",
  1412 => x"1ee0c01e",
  1413 => x"dbff4975",
  1414 => x"86c887cb",
  1415 => x"b7c04c70",
  1416 => x"d4c106ac",
  1417 => x"c0857487",
  1418 => x"897449e0",
  1419 => x"ddc14b75",
  1420 => x"fe714ad4",
  1421 => x"c287f1e9",
  1422 => x"66e8c085",
  1423 => x"c080c148",
  1424 => x"c058a6ec",
  1425 => x"c14966ec",
  1426 => x"02a97081",
  1427 => x"d887c8c0",
  1428 => x"78c048a6",
  1429 => x"d887c5c0",
  1430 => x"78c148a6",
  1431 => x"c21e66d8",
  1432 => x"e0c049a4",
  1433 => x"70887148",
  1434 => x"49751e49",
  1435 => x"87f5d9ff",
  1436 => x"b7c086c8",
  1437 => x"c0ff01a8",
  1438 => x"66e8c087",
  1439 => x"87d1c002",
  1440 => x"81c9496e",
  1441 => x"5166e8c0",
  1442 => x"c5c1486e",
  1443 => x"ccc078f3",
  1444 => x"c9496e87",
  1445 => x"6e51c281",
  1446 => x"e7c6c148",
  1447 => x"c07ec178",
  1448 => x"d8ff87c6",
  1449 => x"4c7087eb",
  1450 => x"f5c0026e",
  1451 => x"4866c887",
  1452 => x"04a866c4",
  1453 => x"c887cbc0",
  1454 => x"80c14866",
  1455 => x"c058a6cc",
  1456 => x"66c487e0",
  1457 => x"c888c148",
  1458 => x"d5c058a6",
  1459 => x"acc6c187",
  1460 => x"87c8c005",
  1461 => x"c14866cc",
  1462 => x"58a6d080",
  1463 => x"87f1d7ff",
  1464 => x"66d04c70",
  1465 => x"d480c148",
  1466 => x"9c7458a6",
  1467 => x"87cbc002",
  1468 => x"c14866c8",
  1469 => x"04a866c8",
  1470 => x"ff87f5f2",
  1471 => x"c887c9d7",
  1472 => x"a8c74866",
  1473 => x"87e5c003",
  1474 => x"48f0f3c2",
  1475 => x"66c878c0",
  1476 => x"c191cb49",
  1477 => x"c48166c0",
  1478 => x"4a6a4aa1",
  1479 => x"c87952c0",
  1480 => x"80c14866",
  1481 => x"c758a6cc",
  1482 => x"dbff04a8",
  1483 => x"8ed0ff87",
  1484 => x"87e9deff",
  1485 => x"64616f4c",
  1486 => x"74655320",
  1487 => x"676e6974",
  1488 => x"00812073",
  1489 => x"65766153",
  1490 => x"74655320",
  1491 => x"676e6974",
  1492 => x"00812073",
  1493 => x"1e00203a",
  1494 => x"4b711e73",
  1495 => x"87c6029b",
  1496 => x"48ecf3c2",
  1497 => x"1ec778c0",
  1498 => x"bfecf3c2",
  1499 => x"e2c11e49",
  1500 => x"f3c21edc",
  1501 => x"ec49bfe8",
  1502 => x"86cc87d1",
  1503 => x"bfe8f3c2",
  1504 => x"87c7e749",
  1505 => x"c8029b73",
  1506 => x"dce2c187",
  1507 => x"c7e7c049",
  1508 => x"ccddff87",
  1509 => x"1e731e87",
  1510 => x"dfc14bc0",
  1511 => x"c6c149c0",
  1512 => x"e3c287c2",
  1513 => x"50c048c9",
  1514 => x"bfffe3c1",
  1515 => x"cfffc049",
  1516 => x"05987087",
  1517 => x"dfc187c4",
  1518 => x"48734bcf",
  1519 => x"87e1dcff",
  1520 => x"30304b42",
  1521 => x"204d3131",
  1522 => x"43202020",
  1523 => x"52004746",
  1524 => x"6c204d4f",
  1525 => x"6964616f",
  1526 => x"6620676e",
  1527 => x"656c6961",
  1528 => x"c81e0064",
  1529 => x"49c187cb",
  1530 => x"fe87ecfd",
  1531 => x"7087cceb",
  1532 => x"87cd0298",
  1533 => x"87c9f4fe",
  1534 => x"c4029870",
  1535 => x"c24ac187",
  1536 => x"724ac087",
  1537 => x"87ce059a",
  1538 => x"e0c11ec0",
  1539 => x"f3c049f2",
  1540 => x"86c487fc",
  1541 => x"1ec087fe",
  1542 => x"49fde0c1",
  1543 => x"87eef3c0",
  1544 => x"f0fd1ec0",
  1545 => x"c0497087",
  1546 => x"c487e3f3",
  1547 => x"8ef887c2",
  1548 => x"44534f26",
  1549 => x"69616620",
  1550 => x"2e64656c",
  1551 => x"6f6f4200",
  1552 => x"676e6974",
  1553 => x"002e2e2e",
  1554 => x"eee8c01e",
  1555 => x"c8f7c087",
  1556 => x"2687f687",
  1557 => x"f3c21e4f",
  1558 => x"78c048ec",
  1559 => x"48e8f3c2",
  1560 => x"fdfd78c0",
  1561 => x"c087e187",
  1562 => x"204f2648",
  1563 => x"20202020",
  1564 => x"20202020",
  1565 => x"20202020",
  1566 => x"74697845",
  1567 => x"20202020",
  1568 => x"20202020",
  1569 => x"20202020",
  1570 => x"20800081",
  1571 => x"20202020",
  1572 => x"20202020",
  1573 => x"42202020",
  1574 => x"006b6361",
  1575 => x"00001123",
  1576 => x"00002d01",
  1577 => x"23000000",
  1578 => x"1f000011",
  1579 => x"0000002d",
  1580 => x"11230000",
  1581 => x"2d3d0000",
  1582 => x"00000000",
  1583 => x"00112300",
  1584 => x"002d5b00",
  1585 => x"00000000",
  1586 => x"00001123",
  1587 => x"00002d79",
  1588 => x"23000000",
  1589 => x"97000011",
  1590 => x"0000002d",
  1591 => x"11230000",
  1592 => x"2db50000",
  1593 => x"00000000",
  1594 => x"00112300",
  1595 => x"00000000",
  1596 => x"00000000",
  1597 => x"000011b8",
  1598 => x"00000000",
  1599 => x"03000000",
  1600 => x"42000019",
  1601 => x"3130304b",
  1602 => x"20204d31",
  1603 => x"4f522020",
  1604 => x"6f4c004d",
  1605 => x"2a206461",
  1606 => x"fe1e002e",
  1607 => x"78c048f0",
  1608 => x"097909cd",
  1609 => x"1e1e4f26",
  1610 => x"7ebff0fe",
  1611 => x"4f262648",
  1612 => x"48f0fe1e",
  1613 => x"4f2678c1",
  1614 => x"48f0fe1e",
  1615 => x"4f2678c0",
  1616 => x"c04a711e",
  1617 => x"4f265252",
  1618 => x"5c5b5e0e",
  1619 => x"86f40e5d",
  1620 => x"6d974d71",
  1621 => x"4ca5c17e",
  1622 => x"c8486c97",
  1623 => x"486e58a6",
  1624 => x"05a866c4",
  1625 => x"48ff87c5",
  1626 => x"ff87e6c0",
  1627 => x"a5c287ca",
  1628 => x"4b6c9749",
  1629 => x"974ba371",
  1630 => x"6c974b6b",
  1631 => x"c1486e7e",
  1632 => x"58a6c880",
  1633 => x"a6cc98c7",
  1634 => x"7c977058",
  1635 => x"7387e1fe",
  1636 => x"268ef448",
  1637 => x"264c264d",
  1638 => x"0e4f264b",
  1639 => x"0e5c5b5e",
  1640 => x"4c7186f4",
  1641 => x"c34a66d8",
  1642 => x"a4c29aff",
  1643 => x"496c974b",
  1644 => x"7249a173",
  1645 => x"7e6c9751",
  1646 => x"80c1486e",
  1647 => x"c758a6c8",
  1648 => x"58a6cc98",
  1649 => x"8ef45470",
  1650 => x"1e87caff",
  1651 => x"87e8fd1e",
  1652 => x"494abfe0",
  1653 => x"99c0e0c0",
  1654 => x"7287cb02",
  1655 => x"d3f7c21e",
  1656 => x"87f7fe49",
  1657 => x"fdfc86c4",
  1658 => x"fd7e7087",
  1659 => x"262687c2",
  1660 => x"f7c21e4f",
  1661 => x"c7fd49d3",
  1662 => x"cbe7c187",
  1663 => x"87dafc49",
  1664 => x"2687d9c5",
  1665 => x"5b5e0e4f",
  1666 => x"c20e5d5c",
  1667 => x"4abff2f7",
  1668 => x"bfd9e9c1",
  1669 => x"bc724c49",
  1670 => x"dbfc4d71",
  1671 => x"744bc087",
  1672 => x"0299d049",
  1673 => x"497587d5",
  1674 => x"1e7199d0",
  1675 => x"efc11ec0",
  1676 => x"82734aeb",
  1677 => x"e4c04912",
  1678 => x"c186c887",
  1679 => x"c8832d2c",
  1680 => x"daff04ab",
  1681 => x"87e8fb87",
  1682 => x"48d9e9c1",
  1683 => x"bff2f7c2",
  1684 => x"264d2678",
  1685 => x"264b264c",
  1686 => x"0000004f",
  1687 => x"d0ff1e00",
  1688 => x"78e1c848",
  1689 => x"c548d4ff",
  1690 => x"0266c478",
  1691 => x"e0c387c3",
  1692 => x"0266c878",
  1693 => x"d4ff87c6",
  1694 => x"78f0c348",
  1695 => x"7148d4ff",
  1696 => x"48d0ff78",
  1697 => x"c078e1c8",
  1698 => x"4f2678e0",
  1699 => x"5c5b5e0e",
  1700 => x"c24c710e",
  1701 => x"fa49d3f7",
  1702 => x"4a7087ee",
  1703 => x"04aab7c0",
  1704 => x"c387e3c2",
  1705 => x"c905aae0",
  1706 => x"cfedc187",
  1707 => x"c278c148",
  1708 => x"f0c387d4",
  1709 => x"87c905aa",
  1710 => x"48cbedc1",
  1711 => x"f5c178c1",
  1712 => x"cfedc187",
  1713 => x"87c702bf",
  1714 => x"c0c24b72",
  1715 => x"7287c2b3",
  1716 => x"059c744b",
  1717 => x"edc187d1",
  1718 => x"c11ebfcb",
  1719 => x"1ebfcfed",
  1720 => x"f8fd4972",
  1721 => x"c186c887",
  1722 => x"02bfcbed",
  1723 => x"7387e0c0",
  1724 => x"29b7c449",
  1725 => x"ebeec191",
  1726 => x"cf4a7381",
  1727 => x"c192c29a",
  1728 => x"70307248",
  1729 => x"72baff4a",
  1730 => x"70986948",
  1731 => x"7387db79",
  1732 => x"29b7c449",
  1733 => x"ebeec191",
  1734 => x"cf4a7381",
  1735 => x"c392c29a",
  1736 => x"70307248",
  1737 => x"b069484a",
  1738 => x"edc17970",
  1739 => x"78c048cf",
  1740 => x"48cbedc1",
  1741 => x"f7c278c0",
  1742 => x"cbf849d3",
  1743 => x"c04a7087",
  1744 => x"fd03aab7",
  1745 => x"48c087dd",
  1746 => x"0087c8fc",
  1747 => x"00000000",
  1748 => x"1e000000",
  1749 => x"fc494a71",
  1750 => x"4f2687f2",
  1751 => x"724ac01e",
  1752 => x"c191c449",
  1753 => x"c081ebee",
  1754 => x"d082c179",
  1755 => x"ee04aab7",
  1756 => x"0e4f2687",
  1757 => x"5d5c5b5e",
  1758 => x"f64d710e",
  1759 => x"4a7587fa",
  1760 => x"922ab7c4",
  1761 => x"82ebeec1",
  1762 => x"9ccf4c75",
  1763 => x"496a94c2",
  1764 => x"c32b744b",
  1765 => x"7448c29b",
  1766 => x"ff4c7030",
  1767 => x"714874bc",
  1768 => x"f67a7098",
  1769 => x"487387ca",
  1770 => x"0087e6fa",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"16000000",
  1787 => x"2e25261e",
  1788 => x"1e3e3d36",
  1789 => x"c848d0ff",
  1790 => x"487178e1",
  1791 => x"7808d4ff",
  1792 => x"ff1e4f26",
  1793 => x"e1c848d0",
  1794 => x"ff487178",
  1795 => x"c47808d4",
  1796 => x"d4ff4866",
  1797 => x"4f267808",
  1798 => x"c44a711e",
  1799 => x"721e4966",
  1800 => x"87deff49",
  1801 => x"c048d0ff",
  1802 => x"262678e0",
  1803 => x"4a711e4f",
  1804 => x"03aab7c2",
  1805 => x"c28287c3",
  1806 => x"c482ce87",
  1807 => x"49721e66",
  1808 => x"2687d5ff",
  1809 => x"ff1e4f26",
  1810 => x"ffc34ad4",
  1811 => x"48d0ff7a",
  1812 => x"de78e1c8",
  1813 => x"ddf7c27a",
  1814 => x"48497abf",
  1815 => x"7a7028c8",
  1816 => x"28d04871",
  1817 => x"48717a70",
  1818 => x"7a7028d8",
  1819 => x"c048d0ff",
  1820 => x"4f2678e0",
  1821 => x"5c5b5e0e",
  1822 => x"4c710e5d",
  1823 => x"bfddf7c2",
  1824 => x"2b744b4d",
  1825 => x"c19b66d0",
  1826 => x"ab66d483",
  1827 => x"c087c204",
  1828 => x"d04a744b",
  1829 => x"31724966",
  1830 => x"9975b9ff",
  1831 => x"30724873",
  1832 => x"71484a70",
  1833 => x"e1f7c2b0",
  1834 => x"87dafe58",
  1835 => x"4c264d26",
  1836 => x"4f264b26",
  1837 => x"48d0ff1e",
  1838 => x"7178c9c8",
  1839 => x"08d4ff48",
  1840 => x"1e4f2678",
  1841 => x"eb494a71",
  1842 => x"48d0ff87",
  1843 => x"4f2678c8",
  1844 => x"711e731e",
  1845 => x"edf7c24b",
  1846 => x"87c302bf",
  1847 => x"ff87ebc2",
  1848 => x"c9c848d0",
  1849 => x"c0497378",
  1850 => x"d4ffb1e0",
  1851 => x"c2787148",
  1852 => x"c048e1f7",
  1853 => x"0266c878",
  1854 => x"ffc387c5",
  1855 => x"c087c249",
  1856 => x"e9f7c249",
  1857 => x"0266cc59",
  1858 => x"d5c587c6",
  1859 => x"87c44ad5",
  1860 => x"4affffcf",
  1861 => x"5aedf7c2",
  1862 => x"48edf7c2",
  1863 => x"87c478c1",
  1864 => x"4c264d26",
  1865 => x"4f264b26",
  1866 => x"5c5b5e0e",
  1867 => x"4a710e5d",
  1868 => x"bfe9f7c2",
  1869 => x"029a724c",
  1870 => x"c84987cb",
  1871 => x"c6f3c191",
  1872 => x"c483714b",
  1873 => x"c6f7c187",
  1874 => x"134dc04b",
  1875 => x"c2997449",
  1876 => x"b9bfe5f7",
  1877 => x"7148d4ff",
  1878 => x"2cb7c178",
  1879 => x"adb7c885",
  1880 => x"c287e804",
  1881 => x"48bfe1f7",
  1882 => x"f7c280c8",
  1883 => x"effe58e5",
  1884 => x"1e731e87",
  1885 => x"4a134b71",
  1886 => x"87cb029a",
  1887 => x"e7fe4972",
  1888 => x"9a4a1387",
  1889 => x"fe87f505",
  1890 => x"c21e87da",
  1891 => x"49bfe1f7",
  1892 => x"48e1f7c2",
  1893 => x"c478a1c1",
  1894 => x"03a9b7c0",
  1895 => x"d4ff87db",
  1896 => x"e5f7c248",
  1897 => x"f7c278bf",
  1898 => x"c249bfe1",
  1899 => x"c148e1f7",
  1900 => x"c0c478a1",
  1901 => x"e504a9b7",
  1902 => x"48d0ff87",
  1903 => x"f7c278c8",
  1904 => x"78c048ed",
  1905 => x"00004f26",
  1906 => x"00000000",
  1907 => x"00000000",
  1908 => x"005f5f00",
  1909 => x"03000000",
  1910 => x"03030003",
  1911 => x"7f140000",
  1912 => x"7f7f147f",
  1913 => x"24000014",
  1914 => x"3a6b6b2e",
  1915 => x"6a4c0012",
  1916 => x"566c1836",
  1917 => x"7e300032",
  1918 => x"3a77594f",
  1919 => x"00004068",
  1920 => x"00030704",
  1921 => x"00000000",
  1922 => x"41633e1c",
  1923 => x"00000000",
  1924 => x"1c3e6341",
  1925 => x"2a080000",
  1926 => x"3e1c1c3e",
  1927 => x"0800082a",
  1928 => x"083e3e08",
  1929 => x"00000008",
  1930 => x"0060e080",
  1931 => x"08000000",
  1932 => x"08080808",
  1933 => x"00000008",
  1934 => x"00606000",
  1935 => x"60400000",
  1936 => x"060c1830",
  1937 => x"3e000103",
  1938 => x"7f4d597f",
  1939 => x"0400003e",
  1940 => x"007f7f06",
  1941 => x"42000000",
  1942 => x"4f597163",
  1943 => x"22000046",
  1944 => x"7f494963",
  1945 => x"1c180036",
  1946 => x"7f7f1316",
  1947 => x"27000010",
  1948 => x"7d454567",
  1949 => x"3c000039",
  1950 => x"79494b7e",
  1951 => x"01000030",
  1952 => x"0f797101",
  1953 => x"36000007",
  1954 => x"7f49497f",
  1955 => x"06000036",
  1956 => x"3f69494f",
  1957 => x"0000001e",
  1958 => x"00666600",
  1959 => x"00000000",
  1960 => x"0066e680",
  1961 => x"08000000",
  1962 => x"22141408",
  1963 => x"14000022",
  1964 => x"14141414",
  1965 => x"22000014",
  1966 => x"08141422",
  1967 => x"02000008",
  1968 => x"0f595103",
  1969 => x"7f3e0006",
  1970 => x"1f555d41",
  1971 => x"7e00001e",
  1972 => x"7f09097f",
  1973 => x"7f00007e",
  1974 => x"7f49497f",
  1975 => x"1c000036",
  1976 => x"4141633e",
  1977 => x"7f000041",
  1978 => x"3e63417f",
  1979 => x"7f00001c",
  1980 => x"4149497f",
  1981 => x"7f000041",
  1982 => x"0109097f",
  1983 => x"3e000001",
  1984 => x"7b49417f",
  1985 => x"7f00007a",
  1986 => x"7f08087f",
  1987 => x"0000007f",
  1988 => x"417f7f41",
  1989 => x"20000000",
  1990 => x"7f404060",
  1991 => x"7f7f003f",
  1992 => x"63361c08",
  1993 => x"7f000041",
  1994 => x"4040407f",
  1995 => x"7f7f0040",
  1996 => x"7f060c06",
  1997 => x"7f7f007f",
  1998 => x"7f180c06",
  1999 => x"3e00007f",
  2000 => x"7f41417f",
  2001 => x"7f00003e",
  2002 => x"0f09097f",
  2003 => x"7f3e0006",
  2004 => x"7e7f6141",
  2005 => x"7f000040",
  2006 => x"7f19097f",
  2007 => x"26000066",
  2008 => x"7b594d6f",
  2009 => x"01000032",
  2010 => x"017f7f01",
  2011 => x"3f000001",
  2012 => x"7f40407f",
  2013 => x"0f00003f",
  2014 => x"3f70703f",
  2015 => x"7f7f000f",
  2016 => x"7f301830",
  2017 => x"6341007f",
  2018 => x"361c1c36",
  2019 => x"03014163",
  2020 => x"067c7c06",
  2021 => x"71610103",
  2022 => x"43474d59",
  2023 => x"00000041",
  2024 => x"41417f7f",
  2025 => x"03010000",
  2026 => x"30180c06",
  2027 => x"00004060",
  2028 => x"7f7f4141",
  2029 => x"0c080000",
  2030 => x"0c060306",
  2031 => x"80800008",
  2032 => x"80808080",
  2033 => x"00000080",
  2034 => x"04070300",
  2035 => x"20000000",
  2036 => x"7c545474",
  2037 => x"7f000078",
  2038 => x"7c44447f",
  2039 => x"38000038",
  2040 => x"4444447c",
  2041 => x"38000000",
  2042 => x"7f44447c",
  2043 => x"3800007f",
  2044 => x"5c54547c",
  2045 => x"04000018",
  2046 => x"05057f7e",
  2047 => x"18000000",
  2048 => x"fca4a4bc",
  2049 => x"7f00007c",
  2050 => x"7c04047f",
  2051 => x"00000078",
  2052 => x"407d3d00",
  2053 => x"80000000",
  2054 => x"7dfd8080",
  2055 => x"7f000000",
  2056 => x"6c38107f",
  2057 => x"00000044",
  2058 => x"407f3f00",
  2059 => x"7c7c0000",
  2060 => x"7c0c180c",
  2061 => x"7c000078",
  2062 => x"7c04047c",
  2063 => x"38000078",
  2064 => x"7c44447c",
  2065 => x"fc000038",
  2066 => x"3c2424fc",
  2067 => x"18000018",
  2068 => x"fc24243c",
  2069 => x"7c0000fc",
  2070 => x"0c04047c",
  2071 => x"48000008",
  2072 => x"7454545c",
  2073 => x"04000020",
  2074 => x"44447f3f",
  2075 => x"3c000000",
  2076 => x"7c40407c",
  2077 => x"1c00007c",
  2078 => x"3c60603c",
  2079 => x"7c3c001c",
  2080 => x"7c603060",
  2081 => x"6c44003c",
  2082 => x"6c381038",
  2083 => x"1c000044",
  2084 => x"3c60e0bc",
  2085 => x"4400001c",
  2086 => x"4c5c7464",
  2087 => x"08000044",
  2088 => x"41773e08",
  2089 => x"00000041",
  2090 => x"007f7f00",
  2091 => x"41000000",
  2092 => x"083e7741",
  2093 => x"01020008",
  2094 => x"02020301",
  2095 => x"7f7f0001",
  2096 => x"7f7f7f7f",
  2097 => x"0808007f",
  2098 => x"3e3e1c1c",
  2099 => x"7f7f7f7f",
  2100 => x"1c1c3e3e",
  2101 => x"10000808",
  2102 => x"187c7c18",
  2103 => x"10000010",
  2104 => x"307c7c30",
  2105 => x"30100010",
  2106 => x"1e786060",
  2107 => x"66420006",
  2108 => x"663c183c",
  2109 => x"38780042",
  2110 => x"6cc6c26a",
  2111 => x"00600038",
  2112 => x"00006000",
  2113 => x"5e0e0060",
  2114 => x"0e5d5c5b",
  2115 => x"c24c711e",
  2116 => x"4dbffef7",
  2117 => x"1ec04bc0",
  2118 => x"c702ab74",
  2119 => x"48a6c487",
  2120 => x"87c578c0",
  2121 => x"c148a6c4",
  2122 => x"1e66c478",
  2123 => x"dfee4973",
  2124 => x"c086c887",
  2125 => x"efef49e0",
  2126 => x"4aa5c487",
  2127 => x"f0f0496a",
  2128 => x"87c6f187",
  2129 => x"83c185cb",
  2130 => x"04abb7c8",
  2131 => x"2687c7ff",
  2132 => x"4c264d26",
  2133 => x"4f264b26",
  2134 => x"c24a711e",
  2135 => x"c25ac2f8",
  2136 => x"c748c2f8",
  2137 => x"ddfe4978",
  2138 => x"1e4f2687",
  2139 => x"4a711e73",
  2140 => x"03aab7c0",
  2141 => x"d5c287d3",
  2142 => x"c405bff8",
  2143 => x"c24bc187",
  2144 => x"c24bc087",
  2145 => x"c45bfcd5",
  2146 => x"fcd5c287",
  2147 => x"f8d5c25a",
  2148 => x"9ac14abf",
  2149 => x"49a2c0c1",
  2150 => x"c287e8ec",
  2151 => x"49bfe0d5",
  2152 => x"bff8d5c2",
  2153 => x"7148fcb1",
  2154 => x"87e8fe78",
  2155 => x"c44a711e",
  2156 => x"49721e66",
  2157 => x"2687f6e9",
  2158 => x"c21e4f26",
  2159 => x"49bff8d5",
  2160 => x"c287d0e6",
  2161 => x"e848f6f7",
  2162 => x"f7c278bf",
  2163 => x"bfec48f2",
  2164 => x"f6f7c278",
  2165 => x"c3494abf",
  2166 => x"b7c899ff",
  2167 => x"7148722a",
  2168 => x"fef7c2b0",
  2169 => x"0e4f2658",
  2170 => x"5d5c5b5e",
  2171 => x"ff4b710e",
  2172 => x"f7c287c8",
  2173 => x"50c048f1",
  2174 => x"f6e54973",
  2175 => x"4c497087",
  2176 => x"eecb9cc2",
  2177 => x"87f8cd49",
  2178 => x"c24d4970",
  2179 => x"bf97f1f7",
  2180 => x"87e2c105",
  2181 => x"c24966d0",
  2182 => x"99bffaf7",
  2183 => x"d487d605",
  2184 => x"f7c24966",
  2185 => x"0599bff2",
  2186 => x"497387cb",
  2187 => x"7087c4e5",
  2188 => x"c1c10298",
  2189 => x"fe4cc187",
  2190 => x"497587c0",
  2191 => x"7087cdcd",
  2192 => x"87c60298",
  2193 => x"48f1f7c2",
  2194 => x"f7c250c1",
  2195 => x"05bf97f1",
  2196 => x"c287e3c0",
  2197 => x"49bffaf7",
  2198 => x"059966d0",
  2199 => x"c287d6ff",
  2200 => x"49bff2f7",
  2201 => x"059966d4",
  2202 => x"7387caff",
  2203 => x"87c3e449",
  2204 => x"fe059870",
  2205 => x"487487ff",
  2206 => x"0e87d5fb",
  2207 => x"5d5c5b5e",
  2208 => x"c086f80e",
  2209 => x"bfec4c4d",
  2210 => x"48a6c47e",
  2211 => x"bffef7c2",
  2212 => x"1e1ec078",
  2213 => x"fd49f7c1",
  2214 => x"86c887cd",
  2215 => x"c0029870",
  2216 => x"d5c287f3",
  2217 => x"c405bfe0",
  2218 => x"c27ec187",
  2219 => x"c27ec087",
  2220 => x"6e48e0d5",
  2221 => x"1efcca78",
  2222 => x"c90266c4",
  2223 => x"48a6c487",
  2224 => x"78f7d3c2",
  2225 => x"a6c487c7",
  2226 => x"c2d4c248",
  2227 => x"4966c478",
  2228 => x"c487fbc8",
  2229 => x"c01ec186",
  2230 => x"fc49c71e",
  2231 => x"86c887c9",
  2232 => x"cd029870",
  2233 => x"fa49ff87",
  2234 => x"dac187c1",
  2235 => x"87c3e249",
  2236 => x"f7c24dc1",
  2237 => x"02bf97f1",
  2238 => x"cdd787c3",
  2239 => x"f6f7c287",
  2240 => x"d5c24bbf",
  2241 => x"c105bff8",
  2242 => x"d5c287e1",
  2243 => x"c002bfe0",
  2244 => x"a6c487f0",
  2245 => x"c0c0c848",
  2246 => x"e4d5c278",
  2247 => x"bf976e7e",
  2248 => x"c1486e49",
  2249 => x"717e7080",
  2250 => x"7087c8e1",
  2251 => x"87c30298",
  2252 => x"c4b366c4",
  2253 => x"b7c14866",
  2254 => x"58a6c828",
  2255 => x"ff059870",
  2256 => x"fdc387db",
  2257 => x"87ebe049",
  2258 => x"e049fac3",
  2259 => x"497387e5",
  2260 => x"7199ffc3",
  2261 => x"f949c01e",
  2262 => x"497387d2",
  2263 => x"7129b7c8",
  2264 => x"f949c11e",
  2265 => x"86c887c6",
  2266 => x"c287c7c6",
  2267 => x"4bbffaf7",
  2268 => x"87df029b",
  2269 => x"bff4d5c2",
  2270 => x"87d0c849",
  2271 => x"c0059870",
  2272 => x"4bc087c4",
  2273 => x"e0c287d3",
  2274 => x"87f4c749",
  2275 => x"58f8d5c2",
  2276 => x"c287c6c0",
  2277 => x"c048f4d5",
  2278 => x"c2497378",
  2279 => x"cfc00599",
  2280 => x"49ebc387",
  2281 => x"87cbdfff",
  2282 => x"99c24970",
  2283 => x"87c2c002",
  2284 => x"49734cfb",
  2285 => x"c00599c1",
  2286 => x"f4c387cf",
  2287 => x"f2deff49",
  2288 => x"c2497087",
  2289 => x"c2c00299",
  2290 => x"734cfa87",
  2291 => x"0599c849",
  2292 => x"c387cfc0",
  2293 => x"deff49f5",
  2294 => x"497087d9",
  2295 => x"c00299c2",
  2296 => x"f8c287d6",
  2297 => x"c002bfc2",
  2298 => x"c14887ca",
  2299 => x"c6f8c288",
  2300 => x"87c2c058",
  2301 => x"4dc14cff",
  2302 => x"99c44973",
  2303 => x"87cfc005",
  2304 => x"ff49f2c3",
  2305 => x"7087ecdd",
  2306 => x"0299c249",
  2307 => x"c287dcc0",
  2308 => x"7ebfc2f8",
  2309 => x"a8b7c748",
  2310 => x"87cbc003",
  2311 => x"80c1486e",
  2312 => x"58c6f8c2",
  2313 => x"fe87c2c0",
  2314 => x"c34dc14c",
  2315 => x"ddff49fd",
  2316 => x"497087c1",
  2317 => x"c00299c2",
  2318 => x"f8c287d5",
  2319 => x"c002bfc2",
  2320 => x"f8c287c9",
  2321 => x"78c048c2",
  2322 => x"fd87c2c0",
  2323 => x"c34dc14c",
  2324 => x"dcff49fa",
  2325 => x"497087dd",
  2326 => x"c00299c2",
  2327 => x"f8c287d9",
  2328 => x"c748bfc2",
  2329 => x"c003a8b7",
  2330 => x"f8c287c9",
  2331 => x"78c748c2",
  2332 => x"fc87c2c0",
  2333 => x"c04dc14c",
  2334 => x"c003acb7",
  2335 => x"66c487d5",
  2336 => x"80d8c148",
  2337 => x"bf6e7e70",
  2338 => x"87c7c002",
  2339 => x"744bbf6e",
  2340 => x"c00f7349",
  2341 => x"1ef0c31e",
  2342 => x"f549dac1",
  2343 => x"86c887c9",
  2344 => x"c0029870",
  2345 => x"f8c287d9",
  2346 => x"6e7ebfc2",
  2347 => x"c491cb49",
  2348 => x"82714a66",
  2349 => x"c6c0026a",
  2350 => x"6e4b6a87",
  2351 => x"750f7349",
  2352 => x"c8c0029d",
  2353 => x"c2f8c287",
  2354 => x"f9f049bf",
  2355 => x"fcd5c287",
  2356 => x"ddc002bf",
  2357 => x"f3c24987",
  2358 => x"02987087",
  2359 => x"c287d3c0",
  2360 => x"49bfc2f8",
  2361 => x"c087dff0",
  2362 => x"87fff149",
  2363 => x"48fcd5c2",
  2364 => x"8ef878c0",
  2365 => x"4a87d9f1",
  2366 => x"656b796f",
  2367 => x"6f207379",
  2368 => x"6f4a006e",
  2369 => x"79656b79",
  2370 => x"666f2073",
  2371 => x"5e0e0066",
  2372 => x"0e5d5c5b",
  2373 => x"c24c711e",
  2374 => x"49bffef7",
  2375 => x"4da1cdc1",
  2376 => x"6981d1c1",
  2377 => x"029c747e",
  2378 => x"a5c487cf",
  2379 => x"c27b744b",
  2380 => x"49bffef7",
  2381 => x"6e87e1f0",
  2382 => x"059c747b",
  2383 => x"4bc087c4",
  2384 => x"4bc187c2",
  2385 => x"e2f04973",
  2386 => x"0266d487",
  2387 => x"c04987c8",
  2388 => x"4a7087ee",
  2389 => x"4ac087c2",
  2390 => x"5ac0d6c2",
  2391 => x"87f0ef26",
  2392 => x"00000000",
  2393 => x"14111258",
  2394 => x"231c1b1d",
  2395 => x"9491595a",
  2396 => x"f4ebf2f5",
  2397 => x"00000000",
  2398 => x"00000000",
  2399 => x"00000000",
  2400 => x"ff4a711e",
  2401 => x"7249bfc8",
  2402 => x"4f2648a1",
  2403 => x"bfc8ff1e",
  2404 => x"c0c0fe89",
  2405 => x"a9c0c0c0",
  2406 => x"c087c401",
  2407 => x"c187c24a",
  2408 => x"2648724a",
  2409 => x"5b5e0e4f",
  2410 => x"710e5d5c",
  2411 => x"4cd4ff4b",
  2412 => x"c04866d0",
  2413 => x"ff49d678",
  2414 => x"c387f8d8",
  2415 => x"496c7cff",
  2416 => x"7199ffc3",
  2417 => x"f0c3494d",
  2418 => x"a9e0c199",
  2419 => x"c387cb05",
  2420 => x"486c7cff",
  2421 => x"66d098c3",
  2422 => x"ffc37808",
  2423 => x"494a6c7c",
  2424 => x"ffc331c8",
  2425 => x"714a6c7c",
  2426 => x"c84972b2",
  2427 => x"7cffc331",
  2428 => x"b2714a6c",
  2429 => x"31c84972",
  2430 => x"6c7cffc3",
  2431 => x"ffb2714a",
  2432 => x"e0c048d0",
  2433 => x"029b7378",
  2434 => x"7b7287c2",
  2435 => x"4d264875",
  2436 => x"4b264c26",
  2437 => x"261e4f26",
  2438 => x"5b5e0e4f",
  2439 => x"86f80e5c",
  2440 => x"a6c81e76",
  2441 => x"87fdfd49",
  2442 => x"4b7086c4",
  2443 => x"a8c2486e",
  2444 => x"87c6c303",
  2445 => x"f0c34a73",
  2446 => x"aad0c19a",
  2447 => x"c187c702",
  2448 => x"c205aae0",
  2449 => x"497387f4",
  2450 => x"c30299c8",
  2451 => x"87c6ff87",
  2452 => x"9cc34c73",
  2453 => x"c105acc2",
  2454 => x"66c487cd",
  2455 => x"7131c949",
  2456 => x"4a66c41e",
  2457 => x"f8c292d4",
  2458 => x"817249c6",
  2459 => x"87ffccfe",
  2460 => x"1e4966c4",
  2461 => x"ff49e3c0",
  2462 => x"d887ddd6",
  2463 => x"f2d5ff49",
  2464 => x"1ec0c887",
  2465 => x"49f6e6c2",
  2466 => x"87cfe9fd",
  2467 => x"c048d0ff",
  2468 => x"e6c278e0",
  2469 => x"66d01ef6",
  2470 => x"c292d44a",
  2471 => x"7249c6f8",
  2472 => x"c7cbfe81",
  2473 => x"c186d087",
  2474 => x"cdc105ac",
  2475 => x"4966c487",
  2476 => x"1e7131c9",
  2477 => x"d44a66c4",
  2478 => x"c6f8c292",
  2479 => x"fe817249",
  2480 => x"c287eccb",
  2481 => x"c81ef6e6",
  2482 => x"92d44a66",
  2483 => x"49c6f8c2",
  2484 => x"c9fe8172",
  2485 => x"66c887d3",
  2486 => x"e3c01e49",
  2487 => x"f7d4ff49",
  2488 => x"ff49d787",
  2489 => x"c887ccd4",
  2490 => x"e6c21ec0",
  2491 => x"e7fd49f6",
  2492 => x"86d087d3",
  2493 => x"c048d0ff",
  2494 => x"8ef878e0",
  2495 => x"0e87d1fc",
  2496 => x"5d5c5b5e",
  2497 => x"4d711e0e",
  2498 => x"d44cd4ff",
  2499 => x"c3487e66",
  2500 => x"c506a8b7",
  2501 => x"c148c087",
  2502 => x"497587e2",
  2503 => x"87e0d9fe",
  2504 => x"66c41e75",
  2505 => x"c293d44b",
  2506 => x"7383c6f8",
  2507 => x"dcc4fe49",
  2508 => x"6b83c887",
  2509 => x"48d0ff4b",
  2510 => x"dd78e1c8",
  2511 => x"c349737c",
  2512 => x"7c7199ff",
  2513 => x"b7c84973",
  2514 => x"99ffc329",
  2515 => x"49737c71",
  2516 => x"c329b7d0",
  2517 => x"7c7199ff",
  2518 => x"b7d84973",
  2519 => x"c07c7129",
  2520 => x"7c7c7c7c",
  2521 => x"7c7c7c7c",
  2522 => x"7c7c7c7c",
  2523 => x"c478e0c0",
  2524 => x"49dc1e66",
  2525 => x"87e0d2ff",
  2526 => x"487386c8",
  2527 => x"87cefa26",
  2528 => x"5c5b5e0e",
  2529 => x"711e0e5d",
  2530 => x"4bd4ff7e",
  2531 => x"f8c21e6e",
  2532 => x"c2fe49ee",
  2533 => x"86c487f7",
  2534 => x"029d4d70",
  2535 => x"c287c3c3",
  2536 => x"4cbff6f8",
  2537 => x"d7fe496e",
  2538 => x"d0ff87d6",
  2539 => x"78c5c848",
  2540 => x"c07bd6c1",
  2541 => x"c17b154a",
  2542 => x"b7e0c082",
  2543 => x"87f504aa",
  2544 => x"c448d0ff",
  2545 => x"78c5c878",
  2546 => x"c17bd3c1",
  2547 => x"7478c47b",
  2548 => x"fcc1029c",
  2549 => x"f6e6c287",
  2550 => x"4dc0c87e",
  2551 => x"acb7c08c",
  2552 => x"c887c603",
  2553 => x"c04da4c0",
  2554 => x"e7f3c24c",
  2555 => x"d049bf97",
  2556 => x"87d20299",
  2557 => x"f8c21ec0",
  2558 => x"c4fe49ee",
  2559 => x"86c487eb",
  2560 => x"c04a4970",
  2561 => x"e6c287ef",
  2562 => x"f8c21ef6",
  2563 => x"c4fe49ee",
  2564 => x"86c487d7",
  2565 => x"ff4a4970",
  2566 => x"c5c848d0",
  2567 => x"7bd4c178",
  2568 => x"7bbf976e",
  2569 => x"80c1486e",
  2570 => x"8dc17e70",
  2571 => x"87f0ff05",
  2572 => x"c448d0ff",
  2573 => x"059a7278",
  2574 => x"48c087c5",
  2575 => x"c187e5c0",
  2576 => x"eef8c21e",
  2577 => x"ffc1fe49",
  2578 => x"7486c487",
  2579 => x"c4fe059c",
  2580 => x"48d0ff87",
  2581 => x"c178c5c8",
  2582 => x"7bc07bd3",
  2583 => x"48c178c4",
  2584 => x"48c087c2",
  2585 => x"264d2626",
  2586 => x"264b264c",
  2587 => x"5b5e0e4f",
  2588 => x"4b710e5c",
  2589 => x"c00266cc",
  2590 => x"c04c87e7",
  2591 => x"c0028cf0",
  2592 => x"4a7487e6",
  2593 => x"df028ac1",
  2594 => x"db028a87",
  2595 => x"d7028a87",
  2596 => x"8ae0c087",
  2597 => x"87e2c002",
  2598 => x"c0028ac1",
  2599 => x"e5c087e3",
  2600 => x"fb497387",
  2601 => x"87de87da",
  2602 => x"49c01e74",
  2603 => x"7487d0f9",
  2604 => x"f949731e",
  2605 => x"86c887c9",
  2606 => x"497387cc",
  2607 => x"c587e5c1",
  2608 => x"c2497387",
  2609 => x"defe87d1",
  2610 => x"c21e0087",
  2611 => x"49bfcce6",
  2612 => x"e6c2b9c1",
  2613 => x"d4ff59d0",
  2614 => x"78ffc348",
  2615 => x"c848d0ff",
  2616 => x"d4ff78e1",
  2617 => x"c478c148",
  2618 => x"ff787131",
  2619 => x"e0c048d0",
  2620 => x"1e4f2678",
  2621 => x"a2c44a71",
  2622 => x"ddf7c249",
  2623 => x"69786a48",
  2624 => x"c2b9c149",
  2625 => x"ff59d0e6",
  2626 => x"ccff87c0",
  2627 => x"48c187f8",
  2628 => x"711e4f26",
  2629 => x"49a2c44a",
  2630 => x"bfddf7c2",
  2631 => x"cce6c27a",
  2632 => x"4f2679bf",
  2633 => x"1e4a711e",
  2634 => x"49eef8c2",
  2635 => x"87ddfcfd",
  2636 => x"987086c4",
  2637 => x"c287dc02",
  2638 => x"c21ef6e6",
  2639 => x"fd49eef8",
  2640 => x"c487e6ff",
  2641 => x"02987086",
  2642 => x"e6c287c9",
  2643 => x"e2fe49f6",
  2644 => x"c087c287",
  2645 => x"1e4f2648",
  2646 => x"c21e4a71",
  2647 => x"fd49eef8",
  2648 => x"c487eafb",
  2649 => x"02987086",
  2650 => x"e6c287de",
  2651 => x"e1fe49f6",
  2652 => x"f6e6c287",
  2653 => x"eef8c21e",
  2654 => x"effffd49",
  2655 => x"7086c487",
  2656 => x"87c40298",
  2657 => x"87c248c1",
  2658 => x"4f2648c0",
  2659 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
