library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"fca4a4bc",
     1 => x"7f00007c",
     2 => x"7c04047f",
     3 => x"00000078",
     4 => x"407d3d00",
     5 => x"80000000",
     6 => x"7dfd8080",
     7 => x"7f000000",
     8 => x"6c38107f",
     9 => x"00000044",
    10 => x"407f3f00",
    11 => x"7c7c0000",
    12 => x"7c0c180c",
    13 => x"7c000078",
    14 => x"7c04047c",
    15 => x"38000078",
    16 => x"7c44447c",
    17 => x"fc000038",
    18 => x"3c2424fc",
    19 => x"18000018",
    20 => x"fc24243c",
    21 => x"7c0000fc",
    22 => x"0c04047c",
    23 => x"48000008",
    24 => x"7454545c",
    25 => x"04000020",
    26 => x"44447f3f",
    27 => x"3c000000",
    28 => x"7c40407c",
    29 => x"1c00007c",
    30 => x"3c60603c",
    31 => x"7c3c001c",
    32 => x"7c603060",
    33 => x"6c44003c",
    34 => x"6c381038",
    35 => x"1c000044",
    36 => x"3c60e0bc",
    37 => x"4400001c",
    38 => x"4c5c7464",
    39 => x"08000044",
    40 => x"41773e08",
    41 => x"00000041",
    42 => x"007f7f00",
    43 => x"41000000",
    44 => x"083e7741",
    45 => x"01020008",
    46 => x"02020301",
    47 => x"7f7f0001",
    48 => x"7f7f7f7f",
    49 => x"0808007f",
    50 => x"3e3e1c1c",
    51 => x"7f7f7f7f",
    52 => x"1c1c3e3e",
    53 => x"10000808",
    54 => x"187c7c18",
    55 => x"10000010",
    56 => x"307c7c30",
    57 => x"30100010",
    58 => x"1e786060",
    59 => x"66420006",
    60 => x"663c183c",
    61 => x"38780042",
    62 => x"6cc6c26a",
    63 => x"00600038",
    64 => x"00006000",
    65 => x"5e0e0060",
    66 => x"0e5d5c5b",
    67 => x"c24c711e",
    68 => x"4dbffef7",
    69 => x"1ec04bc0",
    70 => x"c702ab74",
    71 => x"48a6c487",
    72 => x"87c578c0",
    73 => x"c148a6c4",
    74 => x"1e66c478",
    75 => x"dfee4973",
    76 => x"c086c887",
    77 => x"efef49e0",
    78 => x"4aa5c487",
    79 => x"f0f0496a",
    80 => x"87c6f187",
    81 => x"83c185cb",
    82 => x"04abb7c8",
    83 => x"2687c7ff",
    84 => x"4c264d26",
    85 => x"4f264b26",
    86 => x"c24a711e",
    87 => x"c25ac2f8",
    88 => x"c748c2f8",
    89 => x"ddfe4978",
    90 => x"1e4f2687",
    91 => x"4a711e73",
    92 => x"03aab7c0",
    93 => x"d5c287d3",
    94 => x"c405bff8",
    95 => x"c24bc187",
    96 => x"c24bc087",
    97 => x"c45bfcd5",
    98 => x"fcd5c287",
    99 => x"f8d5c25a",
   100 => x"9ac14abf",
   101 => x"49a2c0c1",
   102 => x"c287e8ec",
   103 => x"49bfe0d5",
   104 => x"bff8d5c2",
   105 => x"7148fcb1",
   106 => x"87e8fe78",
   107 => x"c44a711e",
   108 => x"49721e66",
   109 => x"2687f6e9",
   110 => x"c21e4f26",
   111 => x"49bff8d5",
   112 => x"c287d0e6",
   113 => x"e848f6f7",
   114 => x"f7c278bf",
   115 => x"bfec48f2",
   116 => x"f6f7c278",
   117 => x"c3494abf",
   118 => x"b7c899ff",
   119 => x"7148722a",
   120 => x"fef7c2b0",
   121 => x"0e4f2658",
   122 => x"5d5c5b5e",
   123 => x"ff4b710e",
   124 => x"f7c287c8",
   125 => x"50c048f1",
   126 => x"f6e54973",
   127 => x"4c497087",
   128 => x"eecb9cc2",
   129 => x"87f8cd49",
   130 => x"c24d4970",
   131 => x"bf97f1f7",
   132 => x"87e2c105",
   133 => x"c24966d0",
   134 => x"99bffaf7",
   135 => x"d487d605",
   136 => x"f7c24966",
   137 => x"0599bff2",
   138 => x"497387cb",
   139 => x"7087c4e5",
   140 => x"c1c10298",
   141 => x"fe4cc187",
   142 => x"497587c0",
   143 => x"7087cdcd",
   144 => x"87c60298",
   145 => x"48f1f7c2",
   146 => x"f7c250c1",
   147 => x"05bf97f1",
   148 => x"c287e3c0",
   149 => x"49bffaf7",
   150 => x"059966d0",
   151 => x"c287d6ff",
   152 => x"49bff2f7",
   153 => x"059966d4",
   154 => x"7387caff",
   155 => x"87c3e449",
   156 => x"fe059870",
   157 => x"487487ff",
   158 => x"0e87d5fb",
   159 => x"5d5c5b5e",
   160 => x"c086f80e",
   161 => x"bfec4c4d",
   162 => x"48a6c47e",
   163 => x"bffef7c2",
   164 => x"1e1ec078",
   165 => x"fd49f7c1",
   166 => x"86c887cd",
   167 => x"c0029870",
   168 => x"d5c287f3",
   169 => x"c405bfe0",
   170 => x"c27ec187",
   171 => x"c27ec087",
   172 => x"6e48e0d5",
   173 => x"1efcca78",
   174 => x"c90266c4",
   175 => x"48a6c487",
   176 => x"78f7d3c2",
   177 => x"a6c487c7",
   178 => x"c2d4c248",
   179 => x"4966c478",
   180 => x"c487fbc8",
   181 => x"c01ec186",
   182 => x"fc49c71e",
   183 => x"86c887c9",
   184 => x"cd029870",
   185 => x"fa49ff87",
   186 => x"dac187c1",
   187 => x"87c3e249",
   188 => x"f7c24dc1",
   189 => x"02bf97f1",
   190 => x"cdd787c3",
   191 => x"f6f7c287",
   192 => x"d5c24bbf",
   193 => x"c105bff8",
   194 => x"d5c287e1",
   195 => x"c002bfe0",
   196 => x"a6c487f0",
   197 => x"c0c0c848",
   198 => x"e4d5c278",
   199 => x"bf976e7e",
   200 => x"c1486e49",
   201 => x"717e7080",
   202 => x"7087c8e1",
   203 => x"87c30298",
   204 => x"c4b366c4",
   205 => x"b7c14866",
   206 => x"58a6c828",
   207 => x"ff059870",
   208 => x"fdc387db",
   209 => x"87ebe049",
   210 => x"e049fac3",
   211 => x"497387e5",
   212 => x"7199ffc3",
   213 => x"f949c01e",
   214 => x"497387d2",
   215 => x"7129b7c8",
   216 => x"f949c11e",
   217 => x"86c887c6",
   218 => x"c287c7c6",
   219 => x"4bbffaf7",
   220 => x"87df029b",
   221 => x"bff4d5c2",
   222 => x"87d0c849",
   223 => x"c0059870",
   224 => x"4bc087c4",
   225 => x"e0c287d3",
   226 => x"87f4c749",
   227 => x"58f8d5c2",
   228 => x"c287c6c0",
   229 => x"c048f4d5",
   230 => x"c2497378",
   231 => x"cfc00599",
   232 => x"49ebc387",
   233 => x"87cbdfff",
   234 => x"99c24970",
   235 => x"87c2c002",
   236 => x"49734cfb",
   237 => x"c00599c1",
   238 => x"f4c387cf",
   239 => x"f2deff49",
   240 => x"c2497087",
   241 => x"c2c00299",
   242 => x"734cfa87",
   243 => x"0599c849",
   244 => x"c387cfc0",
   245 => x"deff49f5",
   246 => x"497087d9",
   247 => x"c00299c2",
   248 => x"f8c287d6",
   249 => x"c002bfc2",
   250 => x"c14887ca",
   251 => x"c6f8c288",
   252 => x"87c2c058",
   253 => x"4dc14cff",
   254 => x"99c44973",
   255 => x"87cfc005",
   256 => x"ff49f2c3",
   257 => x"7087ecdd",
   258 => x"0299c249",
   259 => x"c287dcc0",
   260 => x"7ebfc2f8",
   261 => x"a8b7c748",
   262 => x"87cbc003",
   263 => x"80c1486e",
   264 => x"58c6f8c2",
   265 => x"fe87c2c0",
   266 => x"c34dc14c",
   267 => x"ddff49fd",
   268 => x"497087c1",
   269 => x"c00299c2",
   270 => x"f8c287d5",
   271 => x"c002bfc2",
   272 => x"f8c287c9",
   273 => x"78c048c2",
   274 => x"fd87c2c0",
   275 => x"c34dc14c",
   276 => x"dcff49fa",
   277 => x"497087dd",
   278 => x"c00299c2",
   279 => x"f8c287d9",
   280 => x"c748bfc2",
   281 => x"c003a8b7",
   282 => x"f8c287c9",
   283 => x"78c748c2",
   284 => x"fc87c2c0",
   285 => x"c04dc14c",
   286 => x"c003acb7",
   287 => x"66c487d5",
   288 => x"80d8c148",
   289 => x"bf6e7e70",
   290 => x"87c7c002",
   291 => x"744bbf6e",
   292 => x"c00f7349",
   293 => x"1ef0c31e",
   294 => x"f549dac1",
   295 => x"86c887c9",
   296 => x"c0029870",
   297 => x"f8c287d9",
   298 => x"6e7ebfc2",
   299 => x"c491cb49",
   300 => x"82714a66",
   301 => x"c6c0026a",
   302 => x"6e4b6a87",
   303 => x"750f7349",
   304 => x"c8c0029d",
   305 => x"c2f8c287",
   306 => x"f9f049bf",
   307 => x"fcd5c287",
   308 => x"ddc002bf",
   309 => x"f3c24987",
   310 => x"02987087",
   311 => x"c287d3c0",
   312 => x"49bfc2f8",
   313 => x"c087dff0",
   314 => x"87fff149",
   315 => x"48fcd5c2",
   316 => x"8ef878c0",
   317 => x"4a87d9f1",
   318 => x"656b796f",
   319 => x"6f207379",
   320 => x"6f4a006e",
   321 => x"79656b79",
   322 => x"666f2073",
   323 => x"5e0e0066",
   324 => x"0e5d5c5b",
   325 => x"c24c711e",
   326 => x"49bffef7",
   327 => x"4da1cdc1",
   328 => x"6981d1c1",
   329 => x"029c747e",
   330 => x"a5c487cf",
   331 => x"c27b744b",
   332 => x"49bffef7",
   333 => x"6e87e1f0",
   334 => x"059c747b",
   335 => x"4bc087c4",
   336 => x"4bc187c2",
   337 => x"e2f04973",
   338 => x"0266d487",
   339 => x"c04987c8",
   340 => x"4a7087ee",
   341 => x"4ac087c2",
   342 => x"5ac0d6c2",
   343 => x"87f0ef26",
   344 => x"00000000",
   345 => x"14111258",
   346 => x"231c1b1d",
   347 => x"9491595a",
   348 => x"f4ebf2f5",
   349 => x"00000000",
   350 => x"00000000",
   351 => x"00000000",
   352 => x"ff4a711e",
   353 => x"7249bfc8",
   354 => x"4f2648a1",
   355 => x"bfc8ff1e",
   356 => x"c0c0fe89",
   357 => x"a9c0c0c0",
   358 => x"c087c401",
   359 => x"c187c24a",
   360 => x"2648724a",
   361 => x"5b5e0e4f",
   362 => x"710e5d5c",
   363 => x"4cd4ff4b",
   364 => x"c04866d0",
   365 => x"ff49d678",
   366 => x"c387f8d8",
   367 => x"496c7cff",
   368 => x"7199ffc3",
   369 => x"f0c3494d",
   370 => x"a9e0c199",
   371 => x"c387cb05",
   372 => x"486c7cff",
   373 => x"66d098c3",
   374 => x"ffc37808",
   375 => x"494a6c7c",
   376 => x"ffc331c8",
   377 => x"714a6c7c",
   378 => x"c84972b2",
   379 => x"7cffc331",
   380 => x"b2714a6c",
   381 => x"31c84972",
   382 => x"6c7cffc3",
   383 => x"ffb2714a",
   384 => x"e0c048d0",
   385 => x"029b7378",
   386 => x"7b7287c2",
   387 => x"4d264875",
   388 => x"4b264c26",
   389 => x"261e4f26",
   390 => x"5b5e0e4f",
   391 => x"86f80e5c",
   392 => x"a6c81e76",
   393 => x"87fdfd49",
   394 => x"4b7086c4",
   395 => x"a8c2486e",
   396 => x"87c6c303",
   397 => x"f0c34a73",
   398 => x"aad0c19a",
   399 => x"c187c702",
   400 => x"c205aae0",
   401 => x"497387f4",
   402 => x"c30299c8",
   403 => x"87c6ff87",
   404 => x"9cc34c73",
   405 => x"c105acc2",
   406 => x"66c487cd",
   407 => x"7131c949",
   408 => x"4a66c41e",
   409 => x"f8c292d4",
   410 => x"817249c6",
   411 => x"87ffccfe",
   412 => x"1e4966c4",
   413 => x"ff49e3c0",
   414 => x"d887ddd6",
   415 => x"f2d5ff49",
   416 => x"1ec0c887",
   417 => x"49f6e6c2",
   418 => x"87cfe9fd",
   419 => x"c048d0ff",
   420 => x"e6c278e0",
   421 => x"66d01ef6",
   422 => x"c292d44a",
   423 => x"7249c6f8",
   424 => x"c7cbfe81",
   425 => x"c186d087",
   426 => x"cdc105ac",
   427 => x"4966c487",
   428 => x"1e7131c9",
   429 => x"d44a66c4",
   430 => x"c6f8c292",
   431 => x"fe817249",
   432 => x"c287eccb",
   433 => x"c81ef6e6",
   434 => x"92d44a66",
   435 => x"49c6f8c2",
   436 => x"c9fe8172",
   437 => x"66c887d3",
   438 => x"e3c01e49",
   439 => x"f7d4ff49",
   440 => x"ff49d787",
   441 => x"c887ccd4",
   442 => x"e6c21ec0",
   443 => x"e7fd49f6",
   444 => x"86d087d3",
   445 => x"c048d0ff",
   446 => x"8ef878e0",
   447 => x"0e87d1fc",
   448 => x"5d5c5b5e",
   449 => x"4d711e0e",
   450 => x"d44cd4ff",
   451 => x"c3487e66",
   452 => x"c506a8b7",
   453 => x"c148c087",
   454 => x"497587e2",
   455 => x"87e0d9fe",
   456 => x"66c41e75",
   457 => x"c293d44b",
   458 => x"7383c6f8",
   459 => x"dcc4fe49",
   460 => x"6b83c887",
   461 => x"48d0ff4b",
   462 => x"dd78e1c8",
   463 => x"c349737c",
   464 => x"7c7199ff",
   465 => x"b7c84973",
   466 => x"99ffc329",
   467 => x"49737c71",
   468 => x"c329b7d0",
   469 => x"7c7199ff",
   470 => x"b7d84973",
   471 => x"c07c7129",
   472 => x"7c7c7c7c",
   473 => x"7c7c7c7c",
   474 => x"7c7c7c7c",
   475 => x"c478e0c0",
   476 => x"49dc1e66",
   477 => x"87e0d2ff",
   478 => x"487386c8",
   479 => x"87cefa26",
   480 => x"5c5b5e0e",
   481 => x"711e0e5d",
   482 => x"4bd4ff7e",
   483 => x"f8c21e6e",
   484 => x"c2fe49ee",
   485 => x"86c487f7",
   486 => x"029d4d70",
   487 => x"c287c3c3",
   488 => x"4cbff6f8",
   489 => x"d7fe496e",
   490 => x"d0ff87d6",
   491 => x"78c5c848",
   492 => x"c07bd6c1",
   493 => x"c17b154a",
   494 => x"b7e0c082",
   495 => x"87f504aa",
   496 => x"c448d0ff",
   497 => x"78c5c878",
   498 => x"c17bd3c1",
   499 => x"7478c47b",
   500 => x"fcc1029c",
   501 => x"f6e6c287",
   502 => x"4dc0c87e",
   503 => x"acb7c08c",
   504 => x"c887c603",
   505 => x"c04da4c0",
   506 => x"e7f3c24c",
   507 => x"d049bf97",
   508 => x"87d20299",
   509 => x"f8c21ec0",
   510 => x"c4fe49ee",
   511 => x"86c487eb",
   512 => x"c04a4970",
   513 => x"e6c287ef",
   514 => x"f8c21ef6",
   515 => x"c4fe49ee",
   516 => x"86c487d7",
   517 => x"ff4a4970",
   518 => x"c5c848d0",
   519 => x"7bd4c178",
   520 => x"7bbf976e",
   521 => x"80c1486e",
   522 => x"8dc17e70",
   523 => x"87f0ff05",
   524 => x"c448d0ff",
   525 => x"059a7278",
   526 => x"48c087c5",
   527 => x"c187e5c0",
   528 => x"eef8c21e",
   529 => x"ffc1fe49",
   530 => x"7486c487",
   531 => x"c4fe059c",
   532 => x"48d0ff87",
   533 => x"c178c5c8",
   534 => x"7bc07bd3",
   535 => x"48c178c4",
   536 => x"48c087c2",
   537 => x"264d2626",
   538 => x"264b264c",
   539 => x"5b5e0e4f",
   540 => x"4b710e5c",
   541 => x"c00266cc",
   542 => x"c04c87e7",
   543 => x"c0028cf0",
   544 => x"4a7487e6",
   545 => x"df028ac1",
   546 => x"db028a87",
   547 => x"d7028a87",
   548 => x"8ae0c087",
   549 => x"87e2c002",
   550 => x"c0028ac1",
   551 => x"e5c087e3",
   552 => x"fb497387",
   553 => x"87de87da",
   554 => x"49c01e74",
   555 => x"7487d0f9",
   556 => x"f949731e",
   557 => x"86c887c9",
   558 => x"497387cc",
   559 => x"c587e5c1",
   560 => x"c2497387",
   561 => x"defe87d1",
   562 => x"c21e0087",
   563 => x"49bfcce6",
   564 => x"e6c2b9c1",
   565 => x"d4ff59d0",
   566 => x"78ffc348",
   567 => x"c848d0ff",
   568 => x"d4ff78e1",
   569 => x"c478c148",
   570 => x"ff787131",
   571 => x"e0c048d0",
   572 => x"1e4f2678",
   573 => x"a2c44a71",
   574 => x"ddf7c249",
   575 => x"69786a48",
   576 => x"c2b9c149",
   577 => x"ff59d0e6",
   578 => x"ccff87c0",
   579 => x"48c187f8",
   580 => x"711e4f26",
   581 => x"49a2c44a",
   582 => x"bfddf7c2",
   583 => x"cce6c27a",
   584 => x"4f2679bf",
   585 => x"1e4a711e",
   586 => x"49eef8c2",
   587 => x"87ddfcfd",
   588 => x"987086c4",
   589 => x"c287dc02",
   590 => x"c21ef6e6",
   591 => x"fd49eef8",
   592 => x"c487e6ff",
   593 => x"02987086",
   594 => x"e6c287c9",
   595 => x"e2fe49f6",
   596 => x"c087c287",
   597 => x"1e4f2648",
   598 => x"c21e4a71",
   599 => x"fd49eef8",
   600 => x"c487eafb",
   601 => x"02987086",
   602 => x"e6c287de",
   603 => x"e1fe49f6",
   604 => x"f6e6c287",
   605 => x"eef8c21e",
   606 => x"effffd49",
   607 => x"7086c487",
   608 => x"87c40298",
   609 => x"87c248c1",
   610 => x"4f2648c0",
   611 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
