
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"fc",x"a4",x"a4",x"bc"),
     1 => (x"7f",x"00",x"00",x"7c"),
     2 => (x"7c",x"04",x"04",x"7f"),
     3 => (x"00",x"00",x"00",x"78"),
     4 => (x"40",x"7d",x"3d",x"00"),
     5 => (x"80",x"00",x"00",x"00"),
     6 => (x"7d",x"fd",x"80",x"80"),
     7 => (x"7f",x"00",x"00",x"00"),
     8 => (x"6c",x"38",x"10",x"7f"),
     9 => (x"00",x"00",x"00",x"44"),
    10 => (x"40",x"7f",x"3f",x"00"),
    11 => (x"7c",x"7c",x"00",x"00"),
    12 => (x"7c",x"0c",x"18",x"0c"),
    13 => (x"7c",x"00",x"00",x"78"),
    14 => (x"7c",x"04",x"04",x"7c"),
    15 => (x"38",x"00",x"00",x"78"),
    16 => (x"7c",x"44",x"44",x"7c"),
    17 => (x"fc",x"00",x"00",x"38"),
    18 => (x"3c",x"24",x"24",x"fc"),
    19 => (x"18",x"00",x"00",x"18"),
    20 => (x"fc",x"24",x"24",x"3c"),
    21 => (x"7c",x"00",x"00",x"fc"),
    22 => (x"0c",x"04",x"04",x"7c"),
    23 => (x"48",x"00",x"00",x"08"),
    24 => (x"74",x"54",x"54",x"5c"),
    25 => (x"04",x"00",x"00",x"20"),
    26 => (x"44",x"44",x"7f",x"3f"),
    27 => (x"3c",x"00",x"00",x"00"),
    28 => (x"7c",x"40",x"40",x"7c"),
    29 => (x"1c",x"00",x"00",x"7c"),
    30 => (x"3c",x"60",x"60",x"3c"),
    31 => (x"7c",x"3c",x"00",x"1c"),
    32 => (x"7c",x"60",x"30",x"60"),
    33 => (x"6c",x"44",x"00",x"3c"),
    34 => (x"6c",x"38",x"10",x"38"),
    35 => (x"1c",x"00",x"00",x"44"),
    36 => (x"3c",x"60",x"e0",x"bc"),
    37 => (x"44",x"00",x"00",x"1c"),
    38 => (x"4c",x"5c",x"74",x"64"),
    39 => (x"08",x"00",x"00",x"44"),
    40 => (x"41",x"77",x"3e",x"08"),
    41 => (x"00",x"00",x"00",x"41"),
    42 => (x"00",x"7f",x"7f",x"00"),
    43 => (x"41",x"00",x"00",x"00"),
    44 => (x"08",x"3e",x"77",x"41"),
    45 => (x"01",x"02",x"00",x"08"),
    46 => (x"02",x"02",x"03",x"01"),
    47 => (x"7f",x"7f",x"00",x"01"),
    48 => (x"7f",x"7f",x"7f",x"7f"),
    49 => (x"08",x"08",x"00",x"7f"),
    50 => (x"3e",x"3e",x"1c",x"1c"),
    51 => (x"7f",x"7f",x"7f",x"7f"),
    52 => (x"1c",x"1c",x"3e",x"3e"),
    53 => (x"10",x"00",x"08",x"08"),
    54 => (x"18",x"7c",x"7c",x"18"),
    55 => (x"10",x"00",x"00",x"10"),
    56 => (x"30",x"7c",x"7c",x"30"),
    57 => (x"30",x"10",x"00",x"10"),
    58 => (x"1e",x"78",x"60",x"60"),
    59 => (x"66",x"42",x"00",x"06"),
    60 => (x"66",x"3c",x"18",x"3c"),
    61 => (x"38",x"78",x"00",x"42"),
    62 => (x"6c",x"c6",x"c2",x"6a"),
    63 => (x"00",x"60",x"00",x"38"),
    64 => (x"00",x"00",x"60",x"00"),
    65 => (x"5e",x"0e",x"00",x"60"),
    66 => (x"0e",x"5d",x"5c",x"5b"),
    67 => (x"c2",x"4c",x"71",x"1e"),
    68 => (x"4d",x"bf",x"fe",x"f7"),
    69 => (x"1e",x"c0",x"4b",x"c0"),
    70 => (x"c7",x"02",x"ab",x"74"),
    71 => (x"48",x"a6",x"c4",x"87"),
    72 => (x"87",x"c5",x"78",x"c0"),
    73 => (x"c1",x"48",x"a6",x"c4"),
    74 => (x"1e",x"66",x"c4",x"78"),
    75 => (x"df",x"ee",x"49",x"73"),
    76 => (x"c0",x"86",x"c8",x"87"),
    77 => (x"ef",x"ef",x"49",x"e0"),
    78 => (x"4a",x"a5",x"c4",x"87"),
    79 => (x"f0",x"f0",x"49",x"6a"),
    80 => (x"87",x"c6",x"f1",x"87"),
    81 => (x"83",x"c1",x"85",x"cb"),
    82 => (x"04",x"ab",x"b7",x"c8"),
    83 => (x"26",x"87",x"c7",x"ff"),
    84 => (x"4c",x"26",x"4d",x"26"),
    85 => (x"4f",x"26",x"4b",x"26"),
    86 => (x"c2",x"4a",x"71",x"1e"),
    87 => (x"c2",x"5a",x"c2",x"f8"),
    88 => (x"c7",x"48",x"c2",x"f8"),
    89 => (x"dd",x"fe",x"49",x"78"),
    90 => (x"1e",x"4f",x"26",x"87"),
    91 => (x"4a",x"71",x"1e",x"73"),
    92 => (x"03",x"aa",x"b7",x"c0"),
    93 => (x"d5",x"c2",x"87",x"d3"),
    94 => (x"c4",x"05",x"bf",x"f8"),
    95 => (x"c2",x"4b",x"c1",x"87"),
    96 => (x"c2",x"4b",x"c0",x"87"),
    97 => (x"c4",x"5b",x"fc",x"d5"),
    98 => (x"fc",x"d5",x"c2",x"87"),
    99 => (x"f8",x"d5",x"c2",x"5a"),
   100 => (x"9a",x"c1",x"4a",x"bf"),
   101 => (x"49",x"a2",x"c0",x"c1"),
   102 => (x"c2",x"87",x"e8",x"ec"),
   103 => (x"49",x"bf",x"e0",x"d5"),
   104 => (x"bf",x"f8",x"d5",x"c2"),
   105 => (x"71",x"48",x"fc",x"b1"),
   106 => (x"87",x"e8",x"fe",x"78"),
   107 => (x"c4",x"4a",x"71",x"1e"),
   108 => (x"49",x"72",x"1e",x"66"),
   109 => (x"26",x"87",x"f6",x"e9"),
   110 => (x"c2",x"1e",x"4f",x"26"),
   111 => (x"49",x"bf",x"f8",x"d5"),
   112 => (x"c2",x"87",x"d0",x"e6"),
   113 => (x"e8",x"48",x"f6",x"f7"),
   114 => (x"f7",x"c2",x"78",x"bf"),
   115 => (x"bf",x"ec",x"48",x"f2"),
   116 => (x"f6",x"f7",x"c2",x"78"),
   117 => (x"c3",x"49",x"4a",x"bf"),
   118 => (x"b7",x"c8",x"99",x"ff"),
   119 => (x"71",x"48",x"72",x"2a"),
   120 => (x"fe",x"f7",x"c2",x"b0"),
   121 => (x"0e",x"4f",x"26",x"58"),
   122 => (x"5d",x"5c",x"5b",x"5e"),
   123 => (x"ff",x"4b",x"71",x"0e"),
   124 => (x"f7",x"c2",x"87",x"c8"),
   125 => (x"50",x"c0",x"48",x"f1"),
   126 => (x"f6",x"e5",x"49",x"73"),
   127 => (x"4c",x"49",x"70",x"87"),
   128 => (x"ee",x"cb",x"9c",x"c2"),
   129 => (x"87",x"f8",x"cd",x"49"),
   130 => (x"c2",x"4d",x"49",x"70"),
   131 => (x"bf",x"97",x"f1",x"f7"),
   132 => (x"87",x"e2",x"c1",x"05"),
   133 => (x"c2",x"49",x"66",x"d0"),
   134 => (x"99",x"bf",x"fa",x"f7"),
   135 => (x"d4",x"87",x"d6",x"05"),
   136 => (x"f7",x"c2",x"49",x"66"),
   137 => (x"05",x"99",x"bf",x"f2"),
   138 => (x"49",x"73",x"87",x"cb"),
   139 => (x"70",x"87",x"c4",x"e5"),
   140 => (x"c1",x"c1",x"02",x"98"),
   141 => (x"fe",x"4c",x"c1",x"87"),
   142 => (x"49",x"75",x"87",x"c0"),
   143 => (x"70",x"87",x"cd",x"cd"),
   144 => (x"87",x"c6",x"02",x"98"),
   145 => (x"48",x"f1",x"f7",x"c2"),
   146 => (x"f7",x"c2",x"50",x"c1"),
   147 => (x"05",x"bf",x"97",x"f1"),
   148 => (x"c2",x"87",x"e3",x"c0"),
   149 => (x"49",x"bf",x"fa",x"f7"),
   150 => (x"05",x"99",x"66",x"d0"),
   151 => (x"c2",x"87",x"d6",x"ff"),
   152 => (x"49",x"bf",x"f2",x"f7"),
   153 => (x"05",x"99",x"66",x"d4"),
   154 => (x"73",x"87",x"ca",x"ff"),
   155 => (x"87",x"c3",x"e4",x"49"),
   156 => (x"fe",x"05",x"98",x"70"),
   157 => (x"48",x"74",x"87",x"ff"),
   158 => (x"0e",x"87",x"d5",x"fb"),
   159 => (x"5d",x"5c",x"5b",x"5e"),
   160 => (x"c0",x"86",x"f8",x"0e"),
   161 => (x"bf",x"ec",x"4c",x"4d"),
   162 => (x"48",x"a6",x"c4",x"7e"),
   163 => (x"bf",x"fe",x"f7",x"c2"),
   164 => (x"1e",x"1e",x"c0",x"78"),
   165 => (x"fd",x"49",x"f7",x"c1"),
   166 => (x"86",x"c8",x"87",x"cd"),
   167 => (x"c0",x"02",x"98",x"70"),
   168 => (x"d5",x"c2",x"87",x"f3"),
   169 => (x"c4",x"05",x"bf",x"e0"),
   170 => (x"c2",x"7e",x"c1",x"87"),
   171 => (x"c2",x"7e",x"c0",x"87"),
   172 => (x"6e",x"48",x"e0",x"d5"),
   173 => (x"1e",x"fc",x"ca",x"78"),
   174 => (x"c9",x"02",x"66",x"c4"),
   175 => (x"48",x"a6",x"c4",x"87"),
   176 => (x"78",x"f7",x"d3",x"c2"),
   177 => (x"a6",x"c4",x"87",x"c7"),
   178 => (x"c2",x"d4",x"c2",x"48"),
   179 => (x"49",x"66",x"c4",x"78"),
   180 => (x"c4",x"87",x"fb",x"c8"),
   181 => (x"c0",x"1e",x"c1",x"86"),
   182 => (x"fc",x"49",x"c7",x"1e"),
   183 => (x"86",x"c8",x"87",x"c9"),
   184 => (x"cd",x"02",x"98",x"70"),
   185 => (x"fa",x"49",x"ff",x"87"),
   186 => (x"da",x"c1",x"87",x"c1"),
   187 => (x"87",x"c3",x"e2",x"49"),
   188 => (x"f7",x"c2",x"4d",x"c1"),
   189 => (x"02",x"bf",x"97",x"f1"),
   190 => (x"cd",x"d7",x"87",x"c3"),
   191 => (x"f6",x"f7",x"c2",x"87"),
   192 => (x"d5",x"c2",x"4b",x"bf"),
   193 => (x"c1",x"05",x"bf",x"f8"),
   194 => (x"d5",x"c2",x"87",x"e1"),
   195 => (x"c0",x"02",x"bf",x"e0"),
   196 => (x"a6",x"c4",x"87",x"f0"),
   197 => (x"c0",x"c0",x"c8",x"48"),
   198 => (x"e4",x"d5",x"c2",x"78"),
   199 => (x"bf",x"97",x"6e",x"7e"),
   200 => (x"c1",x"48",x"6e",x"49"),
   201 => (x"71",x"7e",x"70",x"80"),
   202 => (x"70",x"87",x"c8",x"e1"),
   203 => (x"87",x"c3",x"02",x"98"),
   204 => (x"c4",x"b3",x"66",x"c4"),
   205 => (x"b7",x"c1",x"48",x"66"),
   206 => (x"58",x"a6",x"c8",x"28"),
   207 => (x"ff",x"05",x"98",x"70"),
   208 => (x"fd",x"c3",x"87",x"db"),
   209 => (x"87",x"eb",x"e0",x"49"),
   210 => (x"e0",x"49",x"fa",x"c3"),
   211 => (x"49",x"73",x"87",x"e5"),
   212 => (x"71",x"99",x"ff",x"c3"),
   213 => (x"f9",x"49",x"c0",x"1e"),
   214 => (x"49",x"73",x"87",x"d2"),
   215 => (x"71",x"29",x"b7",x"c8"),
   216 => (x"f9",x"49",x"c1",x"1e"),
   217 => (x"86",x"c8",x"87",x"c6"),
   218 => (x"c2",x"87",x"c7",x"c6"),
   219 => (x"4b",x"bf",x"fa",x"f7"),
   220 => (x"87",x"df",x"02",x"9b"),
   221 => (x"bf",x"f4",x"d5",x"c2"),
   222 => (x"87",x"d0",x"c8",x"49"),
   223 => (x"c0",x"05",x"98",x"70"),
   224 => (x"4b",x"c0",x"87",x"c4"),
   225 => (x"e0",x"c2",x"87",x"d3"),
   226 => (x"87",x"f4",x"c7",x"49"),
   227 => (x"58",x"f8",x"d5",x"c2"),
   228 => (x"c2",x"87",x"c6",x"c0"),
   229 => (x"c0",x"48",x"f4",x"d5"),
   230 => (x"c2",x"49",x"73",x"78"),
   231 => (x"cf",x"c0",x"05",x"99"),
   232 => (x"49",x"eb",x"c3",x"87"),
   233 => (x"87",x"cb",x"df",x"ff"),
   234 => (x"99",x"c2",x"49",x"70"),
   235 => (x"87",x"c2",x"c0",x"02"),
   236 => (x"49",x"73",x"4c",x"fb"),
   237 => (x"c0",x"05",x"99",x"c1"),
   238 => (x"f4",x"c3",x"87",x"cf"),
   239 => (x"f2",x"de",x"ff",x"49"),
   240 => (x"c2",x"49",x"70",x"87"),
   241 => (x"c2",x"c0",x"02",x"99"),
   242 => (x"73",x"4c",x"fa",x"87"),
   243 => (x"05",x"99",x"c8",x"49"),
   244 => (x"c3",x"87",x"cf",x"c0"),
   245 => (x"de",x"ff",x"49",x"f5"),
   246 => (x"49",x"70",x"87",x"d9"),
   247 => (x"c0",x"02",x"99",x"c2"),
   248 => (x"f8",x"c2",x"87",x"d6"),
   249 => (x"c0",x"02",x"bf",x"c2"),
   250 => (x"c1",x"48",x"87",x"ca"),
   251 => (x"c6",x"f8",x"c2",x"88"),
   252 => (x"87",x"c2",x"c0",x"58"),
   253 => (x"4d",x"c1",x"4c",x"ff"),
   254 => (x"99",x"c4",x"49",x"73"),
   255 => (x"87",x"cf",x"c0",x"05"),
   256 => (x"ff",x"49",x"f2",x"c3"),
   257 => (x"70",x"87",x"ec",x"dd"),
   258 => (x"02",x"99",x"c2",x"49"),
   259 => (x"c2",x"87",x"dc",x"c0"),
   260 => (x"7e",x"bf",x"c2",x"f8"),
   261 => (x"a8",x"b7",x"c7",x"48"),
   262 => (x"87",x"cb",x"c0",x"03"),
   263 => (x"80",x"c1",x"48",x"6e"),
   264 => (x"58",x"c6",x"f8",x"c2"),
   265 => (x"fe",x"87",x"c2",x"c0"),
   266 => (x"c3",x"4d",x"c1",x"4c"),
   267 => (x"dd",x"ff",x"49",x"fd"),
   268 => (x"49",x"70",x"87",x"c1"),
   269 => (x"c0",x"02",x"99",x"c2"),
   270 => (x"f8",x"c2",x"87",x"d5"),
   271 => (x"c0",x"02",x"bf",x"c2"),
   272 => (x"f8",x"c2",x"87",x"c9"),
   273 => (x"78",x"c0",x"48",x"c2"),
   274 => (x"fd",x"87",x"c2",x"c0"),
   275 => (x"c3",x"4d",x"c1",x"4c"),
   276 => (x"dc",x"ff",x"49",x"fa"),
   277 => (x"49",x"70",x"87",x"dd"),
   278 => (x"c0",x"02",x"99",x"c2"),
   279 => (x"f8",x"c2",x"87",x"d9"),
   280 => (x"c7",x"48",x"bf",x"c2"),
   281 => (x"c0",x"03",x"a8",x"b7"),
   282 => (x"f8",x"c2",x"87",x"c9"),
   283 => (x"78",x"c7",x"48",x"c2"),
   284 => (x"fc",x"87",x"c2",x"c0"),
   285 => (x"c0",x"4d",x"c1",x"4c"),
   286 => (x"c0",x"03",x"ac",x"b7"),
   287 => (x"66",x"c4",x"87",x"d5"),
   288 => (x"80",x"d8",x"c1",x"48"),
   289 => (x"bf",x"6e",x"7e",x"70"),
   290 => (x"87",x"c7",x"c0",x"02"),
   291 => (x"74",x"4b",x"bf",x"6e"),
   292 => (x"c0",x"0f",x"73",x"49"),
   293 => (x"1e",x"f0",x"c3",x"1e"),
   294 => (x"f5",x"49",x"da",x"c1"),
   295 => (x"86",x"c8",x"87",x"c9"),
   296 => (x"c0",x"02",x"98",x"70"),
   297 => (x"f8",x"c2",x"87",x"d9"),
   298 => (x"6e",x"7e",x"bf",x"c2"),
   299 => (x"c4",x"91",x"cb",x"49"),
   300 => (x"82",x"71",x"4a",x"66"),
   301 => (x"c6",x"c0",x"02",x"6a"),
   302 => (x"6e",x"4b",x"6a",x"87"),
   303 => (x"75",x"0f",x"73",x"49"),
   304 => (x"c8",x"c0",x"02",x"9d"),
   305 => (x"c2",x"f8",x"c2",x"87"),
   306 => (x"f9",x"f0",x"49",x"bf"),
   307 => (x"fc",x"d5",x"c2",x"87"),
   308 => (x"dd",x"c0",x"02",x"bf"),
   309 => (x"f3",x"c2",x"49",x"87"),
   310 => (x"02",x"98",x"70",x"87"),
   311 => (x"c2",x"87",x"d3",x"c0"),
   312 => (x"49",x"bf",x"c2",x"f8"),
   313 => (x"c0",x"87",x"df",x"f0"),
   314 => (x"87",x"ff",x"f1",x"49"),
   315 => (x"48",x"fc",x"d5",x"c2"),
   316 => (x"8e",x"f8",x"78",x"c0"),
   317 => (x"4a",x"87",x"d9",x"f1"),
   318 => (x"65",x"6b",x"79",x"6f"),
   319 => (x"6f",x"20",x"73",x"79"),
   320 => (x"6f",x"4a",x"00",x"6e"),
   321 => (x"79",x"65",x"6b",x"79"),
   322 => (x"66",x"6f",x"20",x"73"),
   323 => (x"5e",x"0e",x"00",x"66"),
   324 => (x"0e",x"5d",x"5c",x"5b"),
   325 => (x"c2",x"4c",x"71",x"1e"),
   326 => (x"49",x"bf",x"fe",x"f7"),
   327 => (x"4d",x"a1",x"cd",x"c1"),
   328 => (x"69",x"81",x"d1",x"c1"),
   329 => (x"02",x"9c",x"74",x"7e"),
   330 => (x"a5",x"c4",x"87",x"cf"),
   331 => (x"c2",x"7b",x"74",x"4b"),
   332 => (x"49",x"bf",x"fe",x"f7"),
   333 => (x"6e",x"87",x"e1",x"f0"),
   334 => (x"05",x"9c",x"74",x"7b"),
   335 => (x"4b",x"c0",x"87",x"c4"),
   336 => (x"4b",x"c1",x"87",x"c2"),
   337 => (x"e2",x"f0",x"49",x"73"),
   338 => (x"02",x"66",x"d4",x"87"),
   339 => (x"c0",x"49",x"87",x"c8"),
   340 => (x"4a",x"70",x"87",x"ee"),
   341 => (x"4a",x"c0",x"87",x"c2"),
   342 => (x"5a",x"c0",x"d6",x"c2"),
   343 => (x"87",x"f0",x"ef",x"26"),
   344 => (x"00",x"00",x"00",x"00"),
   345 => (x"14",x"11",x"12",x"58"),
   346 => (x"23",x"1c",x"1b",x"1d"),
   347 => (x"94",x"91",x"59",x"5a"),
   348 => (x"f4",x"eb",x"f2",x"f5"),
   349 => (x"00",x"00",x"00",x"00"),
   350 => (x"00",x"00",x"00",x"00"),
   351 => (x"00",x"00",x"00",x"00"),
   352 => (x"ff",x"4a",x"71",x"1e"),
   353 => (x"72",x"49",x"bf",x"c8"),
   354 => (x"4f",x"26",x"48",x"a1"),
   355 => (x"bf",x"c8",x"ff",x"1e"),
   356 => (x"c0",x"c0",x"fe",x"89"),
   357 => (x"a9",x"c0",x"c0",x"c0"),
   358 => (x"c0",x"87",x"c4",x"01"),
   359 => (x"c1",x"87",x"c2",x"4a"),
   360 => (x"26",x"48",x"72",x"4a"),
   361 => (x"5b",x"5e",x"0e",x"4f"),
   362 => (x"71",x"0e",x"5d",x"5c"),
   363 => (x"4c",x"d4",x"ff",x"4b"),
   364 => (x"c0",x"48",x"66",x"d0"),
   365 => (x"ff",x"49",x"d6",x"78"),
   366 => (x"c3",x"87",x"f8",x"d8"),
   367 => (x"49",x"6c",x"7c",x"ff"),
   368 => (x"71",x"99",x"ff",x"c3"),
   369 => (x"f0",x"c3",x"49",x"4d"),
   370 => (x"a9",x"e0",x"c1",x"99"),
   371 => (x"c3",x"87",x"cb",x"05"),
   372 => (x"48",x"6c",x"7c",x"ff"),
   373 => (x"66",x"d0",x"98",x"c3"),
   374 => (x"ff",x"c3",x"78",x"08"),
   375 => (x"49",x"4a",x"6c",x"7c"),
   376 => (x"ff",x"c3",x"31",x"c8"),
   377 => (x"71",x"4a",x"6c",x"7c"),
   378 => (x"c8",x"49",x"72",x"b2"),
   379 => (x"7c",x"ff",x"c3",x"31"),
   380 => (x"b2",x"71",x"4a",x"6c"),
   381 => (x"31",x"c8",x"49",x"72"),
   382 => (x"6c",x"7c",x"ff",x"c3"),
   383 => (x"ff",x"b2",x"71",x"4a"),
   384 => (x"e0",x"c0",x"48",x"d0"),
   385 => (x"02",x"9b",x"73",x"78"),
   386 => (x"7b",x"72",x"87",x"c2"),
   387 => (x"4d",x"26",x"48",x"75"),
   388 => (x"4b",x"26",x"4c",x"26"),
   389 => (x"26",x"1e",x"4f",x"26"),
   390 => (x"5b",x"5e",x"0e",x"4f"),
   391 => (x"86",x"f8",x"0e",x"5c"),
   392 => (x"a6",x"c8",x"1e",x"76"),
   393 => (x"87",x"fd",x"fd",x"49"),
   394 => (x"4b",x"70",x"86",x"c4"),
   395 => (x"a8",x"c2",x"48",x"6e"),
   396 => (x"87",x"c6",x"c3",x"03"),
   397 => (x"f0",x"c3",x"4a",x"73"),
   398 => (x"aa",x"d0",x"c1",x"9a"),
   399 => (x"c1",x"87",x"c7",x"02"),
   400 => (x"c2",x"05",x"aa",x"e0"),
   401 => (x"49",x"73",x"87",x"f4"),
   402 => (x"c3",x"02",x"99",x"c8"),
   403 => (x"87",x"c6",x"ff",x"87"),
   404 => (x"9c",x"c3",x"4c",x"73"),
   405 => (x"c1",x"05",x"ac",x"c2"),
   406 => (x"66",x"c4",x"87",x"cd"),
   407 => (x"71",x"31",x"c9",x"49"),
   408 => (x"4a",x"66",x"c4",x"1e"),
   409 => (x"f8",x"c2",x"92",x"d4"),
   410 => (x"81",x"72",x"49",x"c6"),
   411 => (x"87",x"ff",x"cc",x"fe"),
   412 => (x"1e",x"49",x"66",x"c4"),
   413 => (x"ff",x"49",x"e3",x"c0"),
   414 => (x"d8",x"87",x"dd",x"d6"),
   415 => (x"f2",x"d5",x"ff",x"49"),
   416 => (x"1e",x"c0",x"c8",x"87"),
   417 => (x"49",x"f6",x"e6",x"c2"),
   418 => (x"87",x"cf",x"e9",x"fd"),
   419 => (x"c0",x"48",x"d0",x"ff"),
   420 => (x"e6",x"c2",x"78",x"e0"),
   421 => (x"66",x"d0",x"1e",x"f6"),
   422 => (x"c2",x"92",x"d4",x"4a"),
   423 => (x"72",x"49",x"c6",x"f8"),
   424 => (x"c7",x"cb",x"fe",x"81"),
   425 => (x"c1",x"86",x"d0",x"87"),
   426 => (x"cd",x"c1",x"05",x"ac"),
   427 => (x"49",x"66",x"c4",x"87"),
   428 => (x"1e",x"71",x"31",x"c9"),
   429 => (x"d4",x"4a",x"66",x"c4"),
   430 => (x"c6",x"f8",x"c2",x"92"),
   431 => (x"fe",x"81",x"72",x"49"),
   432 => (x"c2",x"87",x"ec",x"cb"),
   433 => (x"c8",x"1e",x"f6",x"e6"),
   434 => (x"92",x"d4",x"4a",x"66"),
   435 => (x"49",x"c6",x"f8",x"c2"),
   436 => (x"c9",x"fe",x"81",x"72"),
   437 => (x"66",x"c8",x"87",x"d3"),
   438 => (x"e3",x"c0",x"1e",x"49"),
   439 => (x"f7",x"d4",x"ff",x"49"),
   440 => (x"ff",x"49",x"d7",x"87"),
   441 => (x"c8",x"87",x"cc",x"d4"),
   442 => (x"e6",x"c2",x"1e",x"c0"),
   443 => (x"e7",x"fd",x"49",x"f6"),
   444 => (x"86",x"d0",x"87",x"d3"),
   445 => (x"c0",x"48",x"d0",x"ff"),
   446 => (x"8e",x"f8",x"78",x"e0"),
   447 => (x"0e",x"87",x"d1",x"fc"),
   448 => (x"5d",x"5c",x"5b",x"5e"),
   449 => (x"4d",x"71",x"1e",x"0e"),
   450 => (x"d4",x"4c",x"d4",x"ff"),
   451 => (x"c3",x"48",x"7e",x"66"),
   452 => (x"c5",x"06",x"a8",x"b7"),
   453 => (x"c1",x"48",x"c0",x"87"),
   454 => (x"49",x"75",x"87",x"e2"),
   455 => (x"87",x"e0",x"d9",x"fe"),
   456 => (x"66",x"c4",x"1e",x"75"),
   457 => (x"c2",x"93",x"d4",x"4b"),
   458 => (x"73",x"83",x"c6",x"f8"),
   459 => (x"dc",x"c4",x"fe",x"49"),
   460 => (x"6b",x"83",x"c8",x"87"),
   461 => (x"48",x"d0",x"ff",x"4b"),
   462 => (x"dd",x"78",x"e1",x"c8"),
   463 => (x"c3",x"49",x"73",x"7c"),
   464 => (x"7c",x"71",x"99",x"ff"),
   465 => (x"b7",x"c8",x"49",x"73"),
   466 => (x"99",x"ff",x"c3",x"29"),
   467 => (x"49",x"73",x"7c",x"71"),
   468 => (x"c3",x"29",x"b7",x"d0"),
   469 => (x"7c",x"71",x"99",x"ff"),
   470 => (x"b7",x"d8",x"49",x"73"),
   471 => (x"c0",x"7c",x"71",x"29"),
   472 => (x"7c",x"7c",x"7c",x"7c"),
   473 => (x"7c",x"7c",x"7c",x"7c"),
   474 => (x"7c",x"7c",x"7c",x"7c"),
   475 => (x"c4",x"78",x"e0",x"c0"),
   476 => (x"49",x"dc",x"1e",x"66"),
   477 => (x"87",x"e0",x"d2",x"ff"),
   478 => (x"48",x"73",x"86",x"c8"),
   479 => (x"87",x"ce",x"fa",x"26"),
   480 => (x"5c",x"5b",x"5e",x"0e"),
   481 => (x"71",x"1e",x"0e",x"5d"),
   482 => (x"4b",x"d4",x"ff",x"7e"),
   483 => (x"f8",x"c2",x"1e",x"6e"),
   484 => (x"c2",x"fe",x"49",x"ee"),
   485 => (x"86",x"c4",x"87",x"f7"),
   486 => (x"02",x"9d",x"4d",x"70"),
   487 => (x"c2",x"87",x"c3",x"c3"),
   488 => (x"4c",x"bf",x"f6",x"f8"),
   489 => (x"d7",x"fe",x"49",x"6e"),
   490 => (x"d0",x"ff",x"87",x"d6"),
   491 => (x"78",x"c5",x"c8",x"48"),
   492 => (x"c0",x"7b",x"d6",x"c1"),
   493 => (x"c1",x"7b",x"15",x"4a"),
   494 => (x"b7",x"e0",x"c0",x"82"),
   495 => (x"87",x"f5",x"04",x"aa"),
   496 => (x"c4",x"48",x"d0",x"ff"),
   497 => (x"78",x"c5",x"c8",x"78"),
   498 => (x"c1",x"7b",x"d3",x"c1"),
   499 => (x"74",x"78",x"c4",x"7b"),
   500 => (x"fc",x"c1",x"02",x"9c"),
   501 => (x"f6",x"e6",x"c2",x"87"),
   502 => (x"4d",x"c0",x"c8",x"7e"),
   503 => (x"ac",x"b7",x"c0",x"8c"),
   504 => (x"c8",x"87",x"c6",x"03"),
   505 => (x"c0",x"4d",x"a4",x"c0"),
   506 => (x"e7",x"f3",x"c2",x"4c"),
   507 => (x"d0",x"49",x"bf",x"97"),
   508 => (x"87",x"d2",x"02",x"99"),
   509 => (x"f8",x"c2",x"1e",x"c0"),
   510 => (x"c4",x"fe",x"49",x"ee"),
   511 => (x"86",x"c4",x"87",x"eb"),
   512 => (x"c0",x"4a",x"49",x"70"),
   513 => (x"e6",x"c2",x"87",x"ef"),
   514 => (x"f8",x"c2",x"1e",x"f6"),
   515 => (x"c4",x"fe",x"49",x"ee"),
   516 => (x"86",x"c4",x"87",x"d7"),
   517 => (x"ff",x"4a",x"49",x"70"),
   518 => (x"c5",x"c8",x"48",x"d0"),
   519 => (x"7b",x"d4",x"c1",x"78"),
   520 => (x"7b",x"bf",x"97",x"6e"),
   521 => (x"80",x"c1",x"48",x"6e"),
   522 => (x"8d",x"c1",x"7e",x"70"),
   523 => (x"87",x"f0",x"ff",x"05"),
   524 => (x"c4",x"48",x"d0",x"ff"),
   525 => (x"05",x"9a",x"72",x"78"),
   526 => (x"48",x"c0",x"87",x"c5"),
   527 => (x"c1",x"87",x"e5",x"c0"),
   528 => (x"ee",x"f8",x"c2",x"1e"),
   529 => (x"ff",x"c1",x"fe",x"49"),
   530 => (x"74",x"86",x"c4",x"87"),
   531 => (x"c4",x"fe",x"05",x"9c"),
   532 => (x"48",x"d0",x"ff",x"87"),
   533 => (x"c1",x"78",x"c5",x"c8"),
   534 => (x"7b",x"c0",x"7b",x"d3"),
   535 => (x"48",x"c1",x"78",x"c4"),
   536 => (x"48",x"c0",x"87",x"c2"),
   537 => (x"26",x"4d",x"26",x"26"),
   538 => (x"26",x"4b",x"26",x"4c"),
   539 => (x"5b",x"5e",x"0e",x"4f"),
   540 => (x"4b",x"71",x"0e",x"5c"),
   541 => (x"c0",x"02",x"66",x"cc"),
   542 => (x"c0",x"4c",x"87",x"e7"),
   543 => (x"c0",x"02",x"8c",x"f0"),
   544 => (x"4a",x"74",x"87",x"e6"),
   545 => (x"df",x"02",x"8a",x"c1"),
   546 => (x"db",x"02",x"8a",x"87"),
   547 => (x"d7",x"02",x"8a",x"87"),
   548 => (x"8a",x"e0",x"c0",x"87"),
   549 => (x"87",x"e2",x"c0",x"02"),
   550 => (x"c0",x"02",x"8a",x"c1"),
   551 => (x"e5",x"c0",x"87",x"e3"),
   552 => (x"fb",x"49",x"73",x"87"),
   553 => (x"87",x"de",x"87",x"da"),
   554 => (x"49",x"c0",x"1e",x"74"),
   555 => (x"74",x"87",x"d0",x"f9"),
   556 => (x"f9",x"49",x"73",x"1e"),
   557 => (x"86",x"c8",x"87",x"c9"),
   558 => (x"49",x"73",x"87",x"cc"),
   559 => (x"c5",x"87",x"e5",x"c1"),
   560 => (x"c2",x"49",x"73",x"87"),
   561 => (x"de",x"fe",x"87",x"d1"),
   562 => (x"c2",x"1e",x"00",x"87"),
   563 => (x"49",x"bf",x"cc",x"e6"),
   564 => (x"e6",x"c2",x"b9",x"c1"),
   565 => (x"d4",x"ff",x"59",x"d0"),
   566 => (x"78",x"ff",x"c3",x"48"),
   567 => (x"c8",x"48",x"d0",x"ff"),
   568 => (x"d4",x"ff",x"78",x"e1"),
   569 => (x"c4",x"78",x"c1",x"48"),
   570 => (x"ff",x"78",x"71",x"31"),
   571 => (x"e0",x"c0",x"48",x"d0"),
   572 => (x"1e",x"4f",x"26",x"78"),
   573 => (x"a2",x"c4",x"4a",x"71"),
   574 => (x"dd",x"f7",x"c2",x"49"),
   575 => (x"69",x"78",x"6a",x"48"),
   576 => (x"c2",x"b9",x"c1",x"49"),
   577 => (x"ff",x"59",x"d0",x"e6"),
   578 => (x"cc",x"ff",x"87",x"c0"),
   579 => (x"48",x"c1",x"87",x"f8"),
   580 => (x"71",x"1e",x"4f",x"26"),
   581 => (x"49",x"a2",x"c4",x"4a"),
   582 => (x"bf",x"dd",x"f7",x"c2"),
   583 => (x"cc",x"e6",x"c2",x"7a"),
   584 => (x"4f",x"26",x"79",x"bf"),
   585 => (x"1e",x"4a",x"71",x"1e"),
   586 => (x"49",x"ee",x"f8",x"c2"),
   587 => (x"87",x"dd",x"fc",x"fd"),
   588 => (x"98",x"70",x"86",x"c4"),
   589 => (x"c2",x"87",x"dc",x"02"),
   590 => (x"c2",x"1e",x"f6",x"e6"),
   591 => (x"fd",x"49",x"ee",x"f8"),
   592 => (x"c4",x"87",x"e6",x"ff"),
   593 => (x"02",x"98",x"70",x"86"),
   594 => (x"e6",x"c2",x"87",x"c9"),
   595 => (x"e2",x"fe",x"49",x"f6"),
   596 => (x"c0",x"87",x"c2",x"87"),
   597 => (x"1e",x"4f",x"26",x"48"),
   598 => (x"c2",x"1e",x"4a",x"71"),
   599 => (x"fd",x"49",x"ee",x"f8"),
   600 => (x"c4",x"87",x"ea",x"fb"),
   601 => (x"02",x"98",x"70",x"86"),
   602 => (x"e6",x"c2",x"87",x"de"),
   603 => (x"e1",x"fe",x"49",x"f6"),
   604 => (x"f6",x"e6",x"c2",x"87"),
   605 => (x"ee",x"f8",x"c2",x"1e"),
   606 => (x"ef",x"ff",x"fd",x"49"),
   607 => (x"70",x"86",x"c4",x"87"),
   608 => (x"87",x"c4",x"02",x"98"),
   609 => (x"87",x"c2",x"48",x"c1"),
   610 => (x"4f",x"26",x"48",x"c0"),
   611 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

